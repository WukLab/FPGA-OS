`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Cf0Ju7tqgNF03PtViRQp1o7vLG7QVtBfFjlobV/0zdRg4EUwlIJOAGqmc3rxXYDFG9re+1ixCKr6
iq17FH1iMg==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
DhXy9d3szCAuy35qcb4n2WZEInv9fUskYN5FrxT5I9mUTaQuwr0z6lO4SaRk2WIiuLuV6huNnGqa
KiOnZ4KCDf9V7NUBQOG4OTWcJLps/oG2brm3tybE2Q01KttM3NytG5iDziOahBTaKwqT+CP5NNcL
76iBNr/u+G2jxi4ludw=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
NUv2qb8xKeaXgyk5a7IPSw6Mvsu+RfDjC1v0WcvyV1Dl5cS8enBwd0FPEGRO3ZBL1Q3ASB/VlbTw
N5nSW3Q/DzR1Ng9qbo7FpUbmBa70IFOrAzJIRGsgzMpzG3j7r8C7rkvjTfU+qjkTC/r5opgqpAqC
hio6UL/OlNYCYRfMCH8+kImjrwhYxx6YVfe2J9TcGYBJ4KKNsp5ONc2Ty+vutRmIkuOa//YeFDM+
xhU76i5YWEXERyItfHjpta06PhPcDxxrLEwkaJlIMrBM0ZBO8NsxGZNeWkOoTPuOYb5am6WqFK+D
r3oorQhZIHrxkXZluUm2QbVHT2nQzfke0ruXKw==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
P5Z29ozOqi1XRTudJDTzEZms1i4PR0a3QiMg+2woopusY4Bgbe6NiumhjvdT0KhoZ2uS2GOVkhLs
Nn7o7HmdYuH6EgdiomHcj3zME+Bqqgfxi5F4HGzxtcai9kWd5tewkGUeMzlfe4xJKEaJzoecxMBk
pgobQJmz34epe+DTY2K0oSl1BntC5yc3wdlgzcDh+xWKk2ivHYBGyZMjE9ByN5eso11iMxaHv2I9
Pi2GiPgyexH8t35GTSBPH8+a1df/PQwvPLAuiYi96JjIzpubTAY+ATuT8VZelBGW7eXHI+OIwSOn
Gn5dCw2EnfCaWoGd1pJD6jATJ5cBIztjLsCFjg==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
BXCYl5tBQ7RRFptBJgUurkZkIKGuDwhxSFIBoNWZxJ3m+klqoerKzegP81LuiinTzQTP1jvpxbUI
m+mbG16pnuceVHdORvZRYH1Vizu1VQTykTI6wUafqjyusX/BtF/P4dJo/NSUW9sjw2yGhlXku9XW
7N+WY3mHvt1cyuTCQWywWBlGnlDJkX7qcHxusY0MkGEsW8P+fyqr87Dj43e0HVrpxyYPcWRitIZk
OcDzPZYt912Mb7xAgBrOVlxHwDAT994giTTN4U9EhMgLI83GOdHN3dbbADqjj3lGZcw7Q0x+MIFj
BRSQALyhmkO2kHexlaIrSA1aYt8PV3+aCwmYIw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
fyVU8xm5NYWN9sEAIlJfL4u/hp6kbCsPQeW9z2eGGl9mL/SsXCxPdevSiV4Bslj1S4o9bDuhzIfs
gKAJfgOvzQjFzu9mluxcXNjHeplTB3jixHgIDEqZwDlCHJvplWcXHilcXd9zstRK5lqdAGTRgydp
3+0Dg7xTJTYPEQgyTaQ=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
T5GlPDh7jS+EYlaA9KS+YN1MT8pan/Z5Ia0YJRRzqEBBafOxLT6fBxc4ej+CZomMShslPQonqHPQ
9cAn0hwj19jZ7k03Q5cvmqHJizeQyCy6ZoDwqqW385Ef2z5Wkc/SFD/3eVNlAo/N5JW74EgWFaUm
U67gl4V5HYtvvbf95mxjf9o6VBtmhgiDnoF/BYmquumejBMSnMqwMXrlZPUC01nbLCucBXNL7xdL
CPgRKL94BD5wrJXndQv8Hfvmvgmzx1cDOirI23QFaaM9puZOESjeBMnicCHPf5pE9r6uswbIjOPU
E92+926TozPYBXCXRaS9wHlWKOA4nXmsFWkQFw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 151824)
`pragma protect data_block
0JnHFdJlY/sagd6Qfal8PBbMoWfeE/GHiFP6ED/4Dcm8eEuvF892DRIDPEJqY6+qYcuIdF9uXpUQ
QZmFcGBvJRiwvoF/GP11xKVjlrU0k4ubSP+1yR6m5HNbPUzWv+eDy+Tm/FaHSUUE+t32Zsiz46Ht
aaf6ECkvyCkeBjZID+XwDgXX82Mu9IFmpknjUVeSYaijCzlm/VEcvn1oP7GJjL01oY71BAOD0/Rt
V8YMZjqczSiyuQX7BYvSmedOK8nX+1hHP5rbaNg+hdK8Nq3YPpRP4RR0/MYhYMofT7O1Jcb9SS5+
awy1pFh4pI3AMpJBQJmxUybdti2UxU6pL6AJPmMQPpGZNF8d+Q2Bx9Ah3uGncrb7UDXdGhEiyvjV
8XHso0qfWedtLKlcGCezw9iC8duNwSv1GJFVyfsTYZ4IsVufJPg5/HcE+eq/kZ0v7/Ofop7TNhrn
N3QSn666I8CraBDN/NYp1ze2NFdIyXQ7OxqXoj4lo/C6+r1YtVMvpOTvGZ+x8xPM8Rf6gBvQ8Y8G
FtIsb40Wv2ldYeFgdHzzF5aGObmioJBZdxoDVqM/GZEvagkK5ET9dAw3Kod2DpJfjf7ok4j2Gays
PCJ8lnf6h737kLQEAN12tIP/wIkWJN2VQyBw+IPSMWkA/tD1Fttm0j4fiNb7q7gqjHBzSw3ph4hd
355yaD2tMEhWst+kDNAsMivEVPKNZNSgn8lZPRFHc50VlNa+Zuhhivz7qTLAVv6WiPVLQTJpdWhh
6DkTa5Ki0qEohNcoEuRvjiZQ+RsIBtmR0jCXqN8Jmj+kDTxE+3ni0hULbSAgaYNObp6cDsVdWprx
dFKqSBG8jQo5t2nUnTU7+Y0rDgbyw0qVBgaoGt2ICtI2k1OW09wgHwG7jTlaUVMVmQUKl3wuWQuJ
sQTZDzmSWscg51kDSUzQ+zemTG/lg1mrgx4xiXRJe8MpD18c6SGamn6q99BX0N7OrzpbtyF5s6x/
QLHzGvv+fPlmWo59RAWE7Vl5iE2iYhXcnm4SXRgIS8HOxz2MGYh1VXJkLlpQBwyO+xTr+I+2shTe
iCIFr0MpnEfHpLUF4Ii3iLq+WeK/h7E5HxKToBJfKdNtREbmITcuQU822AECgY1Cp047XI17ouuu
QutZ5o/jwMggrC4VfrU4xf6WJVob6SWLrs22KI1MJeg9ZfHgoWBKkGmtcCupcLMZfqE3A7GbV8Jl
kcAVWuFR2MBRWo/jnz3QBBkXUTY2vcpidJBoJiMG1HpANz6TvhHqaePKRk/icHomb31ZNBjTjNi1
F+U1t4IAPRQCVKYURWbcF3vf87wLyVL83r65a0sJlH9E9TYxlC/dEhi7Y82KA3eTzEdg6wRKGdkU
0wepcxjlye5t3IojmzmRP5qeah6Y3QFjpA3FAfWvPZHRDya0G3WOkrUmn4TvCqtc6dO+VCSoM7r6
k05SdcSzXi2NKj58Z7zNql3KHHkFBMTmcA02pqCkzuUwuuJa/HAkv+ZLUkR+38cQ+L/mJpUyJHrG
KGXp5tx2WC/K7q2cR7wX0kDWVBTHySMSXjtjB7CnEQZ1aDPZ3muVxLFBujj1uWrpWjHe54DGXT5O
JM2nobmUxf3g8FVpQe9fyuhcbqC85NAglXLTiowxx0C6A8S7W5APTOx8n98WBNj70yGru7n1Ppoq
p0RHnoLUjUSbpd5rQCY7d8ZTA6JGhywruST7MYXQYg29dQM2vbSSA/tsPNrhGU9N6JmYVU/1yvE2
3WsgXq9hXdrbqV5Ihr3QTLVm6oER9I/bVEsDjFFAYPJcurDUTyEVYjdpYcIyeT1DsKwuKGboV19L
bPSPkL0wOryvYQF5tkXf5PHwpIBHnQsJVchlw1ALmRLxIL7tGT9QKxpLIvfng4Tru8zKtI8DnUsw
M6eb4wtPKNlnDOaM4RUfVJeivZdBKySvPmkZuT/SQ91/gzKWzsfjD2uYYtmh4p/+AAzTJEfW9Q/c
EC37HINMqVSvBHezdNIZ0pvcnYAM1ocPkecVLCOpWWsmCmvXnHVQ/yfFr9XqkiwOri9CXxNcJjpg
zcqQ6TT+njJvYHU3dLUKgKMgU9O9E95Eeq0ai3II0EHqWkNrhxJnnEnGp7+wxl3m4zEA0aqsn2/g
v4bADEADUfn1Yz7VqzHOVGAQPvuMFhblhgK4GuZrhVCcSw43OMcSLFPXd2Od34JLRd1W8rRtOiCY
aYkTBnlRPlU9VpsufUVtOaydpVabI43FzGAkPaQJ33yxorZPVms04LmSHRsB7MsI3sFM6U/fRSF6
K5FP7rfWhgOvjTaqmB0j+hDYJMDJiO130JzJgwSMtyGQtQi4GyZFZzomsQyUQvyqTVVGocf4qk9Z
qEHOAfn46h4lJunmfpF/LI8m6BrAB4bkq/hcWLCVlCjfx4Fqe8VGHaJgpj++usECBmqZe7ff6rfS
MQivjfh3ZeyGH5CI1ijSQg+dEEiFR6Qqa68YvUtHFVb2UUSzCwi//bV3VSvAw1hOO2F2ckymlRfv
iPhctRMcFenfIuiTumYMRAa0lAcLhGypkcw6dZSle12APU80Q3DI5FEAdZXRzsBll3er6u9z6AkD
RsP6ZZw4AKL6LOJ0HSbUYy64jsUG49phHEiVtbP8XMnQf795TTB5Uk9QAvelDEbZDb0gG1DOGAbA
oiuvlbhjeNth7cfnwDCrjCrajoGAbD72SBiZsksNEECeWlp/6XIqZcZcybpw+pHvHaMt3nEsAWBY
6Mfp8hEFZPLZOWIuYDknok/0C5VVmBgpngF2vFXeyNfFuScL2K+dghf1Xqd/dCOUyD5QApKY0FFE
U+7MNTrBhjMpTBNYFX76Jy0+7DIfYjsXsbADhvQzzzAw6bdbnEH0AzJHFQSO7Iv13b/yX6pmp81g
xYV4sybR06BRy/2g+qOlllcrG8JdcsfZ8Rqm1PikSsk+Qjb4xKF6Ka1D0MFhIrL+RUhnyq37thsp
ighI0sKQx0Ex8znNqLNzMt3k5hmR0CCi89oyWkfpnV7hiH5I3In8bQeXENZMuhfKkVGIbW+gqkXO
+at4WVG2Z34iTOer2Jw8NvtWjqZKqMI8VqdjRNXk6NrC8S3Gt/u4xVyLYKJiViyWb98Hyvp/hLxi
yXr6Mq07Kf9QdIwHiBezDswcQxzIYZm43Ifdp8tAsHMWIYywKKG7/h375V2YApRgo04n3ry7Psxp
JRGH+Pt5YKXGY/ayhBg3hxh0cGHmH6sRnAtWEBB6ErIwonWIxDCxGxVdWGd6rSQiVUABEpva8yaM
L57sETiUrJNHOrYoDg3dZfaohxss4wYQlsDql80od6Cr1vZq9f7Dz+tby3IBCjfEd226P2B/Qswn
iMZ5QJO4D7T+5+E81gOsa0zd3Vugyd7v8FGiuuQIsQc4rVqDxuAqrTV/IZIFZk2sYwrFhc9lgQMM
HgPjJBsOa9jLN2GeaMz4vDyitZulI6j4Bkk4aXPKbjZlCIOpyXScyhaYEz/MTle+PURW1TEmKJ3I
Neqe8XNcVz7vBChugRo1Eh6dTU8h469TkNnmcZEse/9vyv3AygsHkpKLMWpv3eShc6wZku4lpZwn
v2ubWqxOplwj5+9lSLeMkXaGR2BGUWJlb73x8YEyaezWqU8RIDEhEMlERB/lIfQHoA1v2rfZtOnC
SNWcj8jiXqb8bDoQKwUgbK4inzEjlzJCL43g7i7qgBg/kQCskbsltw/f+nWU0ZJIJpMjpJZkt+yB
zqCYsuQiIdM2ldGO/E1VjvxnLUnWk4U8Nf+Qtaj/RUmepl+m5gkkTmZGAHJPKCXv8Ss9kQtPGKhq
/jXlABqpbPtvvC7FOin0lbcbkieB98mObDCqvhdTO4aTfrMI/HsYNyQoS/okxqLcUUUs9vdmSNWU
4riU47CrAqDatNIls9je4dKxVWmYf83SqIlfP8/Llk+X3IkAHkv3p0s8Vp6fF1CFSkNs3+FKxE9K
fnkigklVyrRyiBJBSciOB65EUAUWWNkGcwfZa66Psd9GOIp9w9yudB9gtqHYiSDZAsC7GuxVuKUR
b+C+qdltZW/Syx4zhK59hxZuLqe/R0aHwwXojBg79fTm2NMh2q2M0MqKgK6OWny9yNHEZAs6Nk04
JBWIOUzK/PfajN2WZCTS0ZnBIE/wWuWZ9yq2r3qntgmOvkdQeowMxwKvB+IWjYG8XIG8yPmiO+Dr
VlFb+CJuITfyPujcB3VpfcZdIQrjaYiQvpdMSCF8tTvFaSdqUEUym2tB40kNhVVRuTxHqvNFesAu
3ydXShN+BQDDrIXVeVoAXloLgaXjxmj5JDsYdedPju88qjDbtrDU5cnSYImg/v5ACNZTAQ8NbFMw
jca9c0BhClzIgY5bl1LLSIF3hxqKeK9rgDk+1+CxkNQVmKzk9GBTakQjZYIiRxPGpZXn+QXG8wZa
AL9DZVl/3yoET7kE4cqhTFb4TmB2HdTSrhkmK/oJxAW14vuUYcj5cxpHDYDWef8VTobogA+LIGZj
hip8sKXTyg2f2vsmKbYbxzRBg2Ufdzb3isPvzeKUN2RHvR4URqKd5KOeRmtwbzj+oBguH1ZubTae
LPB3bA6PGWWEvzBqvkpQIdBmYnx6Iz9OIieEYpvoPtPPXo+7GH/385K1iMy8CBIDEiApV7BuS9Zf
47gPqhVgphnQE1BkuWr06CeclAjV0/3IF4Oe/BAdIuvIWxh35Q3XB+SGIQqt1Ec6WqMmZjb18xvt
kZ/i9+jrXvhfLTSylwCI6aFaYlUJES4EUduzwZgrNCrIULI51aZ58Ej1kc83uzUkR9wTIqRAUpQG
frGTviX1VndkErGFPzCBwcOrsrUZgR3TnddLsjI9Ft7tAt+MB9HU9QVKXu9wMsUZa/d6pSDJe/O4
gH1jM2ExT1gwDvmFOoBtYIvY1Wiq5eg7gON8WiXAETmcMDLiY5sgkpLMv8xe5GXoDpAx39xVzn0v
rr0v4fnguWkB+K8MlFW0faEXc+Npe2L8amwuqki7UvVtT1iZ0dI6/5ZD1ofAnfg9QXS0M9dYur5n
hKYh7lAz6BOnWFsyI48lnvbB5+Ne6VRI582ojsPO4gjAfYm9D+9FIHtzxlOriDzrE+xolWfU4C2b
xFcBNjOlpQjFLX29AWtSrnp4A967zWRpsWSIdslCytsM/T50teIujTxasdePMo6RV8jNM/mXqzZy
6mYDgS/ldtil9dq3PwbRswxXyKDgWEMrh2a/dkAo7UWk+URm+tp/jy7KAJZgYo4oB/vtYR4iWOxB
jOly6YEIEXZIoPPMZrJpjGXLen1Q3mzHbiUNwKe7ueuuJ99T6Rdq9Rv2+iGPl8sQfooU1b4yKFCB
nxFo1icmRd+mTESd82WF8NtYtT7j8oYPJULxxvF7by+lTyO1iSKBBQxISV230FkAaJS+gYPoMDMU
L3UZmJj2TQI1ZifOggrKqcP3mC59ZHL0TOQB98BHfpKE0l4VKTlsxW14ucJe2GOa3DZ2b9W2Sf2P
avCnllnUMCxb+CFxgpzTm0pqV5V+PyvXH4nI5qQhF6jVtbrPqRrVL2RnXtfmNzMxhJeSnJsHHIeL
RyPePaxSR2iTMIacRy9UfIaaeGtEcLIrV0KvPqZaFMNes6VBnv8sfzparxkYLOP1gDPAK//DPjbn
TpEGjmemdx3FGi+j4Q564ZAFsxyPzAE9kDAh3i/57L7I2J+vnQCDG5beBSjqt67eMIImfidPoxhy
QpGA08rCxTEkmyKVcUUmPSSgJfwpfY4t9ExkS1FM3I+P6WeeyUpzWQGOEM9eAxiMGEF228D8a7oT
YVdPXhYOcH2DgudtUcuqgDQ8LssO/TX7H41SO9aQRqOl+C1KbAOsOqleOwNj3Ykqk0H2hs8JlEP3
pry3b7/coHokNyMH4EZC62aJ8WoVObAGuUh3xG85+I+3kMLZaoAr36AXo4R2gyU5uT628Te25fZe
FPO6iL7kBCGPAyGsnnbhsWQCLH62ashXIKev/P3R/hBSU7YnQyrgWBpR1y03f4urLr+em/LQs2WR
+SD15QqZKvXvfWKbN7mUHz9raZNC+an785IN4ohgpfLN3OlWImOqqV4EnwCY0/xLD9AfG4VhjAL4
Yi5dnRMeFN87OKA00N6fVX8CcbA4QCjlUIFF7QbfdAXyjNkoR7D3Zp578RfXPKDg1hNPixDJekBV
NM3NJeWksrxY8aBqTdnSvC8liRnMT1DKcSgg7Qclo0e6WR6t409Y63u3z4u8gzs/faTHD3EUIxx6
WHyK0A4nMyQ3bfTYeg1XTPwDvMqxx2JUaC+KbXyBi8OzVoxCEMZacFtIHD4jUbG1AD+Jsbn7rfVY
Jy5TVtlPbmCpcJnuNQIPUyrUIoyDcG86qmg+yQ0Y9mvz8wMrD67CVxJrie3DaE7CLDhy66NJDJsu
3BejvY0anhr/NhJodxXNzszeUStBGteIQ0UopBYbeOiUtu+hfe7soMi3QIa0GFudJzq+1WmrD99y
de7EEJd84ofLKeXu0REeC2jjBRpu4H235ejM6n2xx26Uxfve+C+gfKsWZhXynFHPyljjgrXjEtRD
4wz50PFpEk9TXFtbM2Rvp1N3ugt0hTLn4swuRl3fxemQqhaPZ2Hoq7tGhoduIy0LQzbfjA41+512
6pDDOQ6+qEVR59osPwvsxvvRMiYmJBM0anqb7daI7bW33GKDpOBxx8t0BiO8nq2fm6MseqZ3QQVI
b3Y0O9TikkT8R1TtffE8Ti5borIa5kY8q9wbm/JJMta9AdqJ0ntxpUTd5OTRy7lw1TH27N7SB07e
KzkgQXBuXr0O+B+ry1ORdLJ5zz4yAWQcNCcIxbpIDNl2xyGHBLiHqJeAUAYngaA/TAe6oNHNd9+t
fue5sSGaro+J2EqCOUOn2yFkFD79u7CJBhXZUCaw+CzQo6FoZ4PKGdOQnORACVp5/2SyO8R5btp0
ops2wvcwuv9ntr8CYg5Rrd+bsxagnjr+bOLvvCsQpe/c75usX8Ur4ey/GleCgyq2bs0yPZJcS9Fw
QhexiB6sqwbjkPCv27zymmgM65oxOAaCtkvFAFwAqeoTCAwpzJpW5eJfMdjQQkwj/of9AhTmH603
8ukJctvWCbM/ftRjvCRHws2cjufVYbaFo3+9Y/B2Y78CqpwqnYcQ0Pt//uw6EOyM7o9+CL8woAr/
0u3RaXYg2iYuNOwggajeo1TK1U+PRVGicmNWaQIdOTZUxjW8+Vt1b73WU9vrr4sM85hc+F4lxEcN
Qp/u0KIh2kFNyYfbgxKQ5z6cCEm2jbtEG5gTVlupSnZwG4jE66NAOqPTZj8cS6XhUDe4s8Zr94jY
PSzS7sy0NCvJMnCASqRt+1jPIPC7CKlHDy2a9TbEkAOZ3AqIShhxMyDKmzOEag48JzIV5V7juyh/
VWX9fTLHcUKcSqAXmqHgmL9zXF9Zt1RkpJNPxzAx3Db7++PaMMq9Ah+Txr3oAHvApUG+q5WVa/XC
MSrcv/3ETU08OvaOPJ/0iHqA8GZd0wyTLsbyaw+8YYyH6xKlz2j/mphB3Pum20jGRLtAC5aEVpcQ
ZK19gOGLlJMx+7Ptlft1VLb2RLsl9pqWJvBu1ykq5P7F8BFTNIjJ4CqqhpR9Flm+lY0ULM/1qiq/
FCUDkGbr6zsrPV6GP+boKrDTvfYljVo1Hgc6pdx+oidAXhgYcRfMsqpKdmpLKmGHwLKkm/GNhP4D
OIsQq+ux80MPTrDK8ovUnBbvD4LeupM6wgXX61bEguRB/G+EkALIQxG7vvK+Ta+omCVAOkMmeLyn
Y/mPu0DeCSxueTBwcHWhyKq/mXfJlhu3U0ab2zKw3TceuwQ9i9nD0BvFefjApqvP4tvOpKQqNC3j
KvXC4Pi7wPSXm5+HfL6cJTqLR1NHSKLS2q6UM6f10QBDlUzpkuN6bmT+1zKrbHl057mAvm0jUwMg
zZIb/vWmq3RvKCPJhG/Sz6h5BAHPm/Pw6/TX9u2dAJbNk7cOGxY/pw4RFjQ2xESfKs6mEJ+UBbjQ
AzPtq3ibwqJObH2zQaOR1xcWHXahz1OvuA4J74mUVSS8Fpphov6t75Uw9h6ooBJQ+m6Ww4aMWqOP
aWZ5P1RqB7O13VbVoxa4xziTP6pcSGwij4cXLFf5xmyfO/ogRdnkkoegGFI1U/R69DzPqQTiUuXn
X4nKG/PAf/1xJOXCRYxNKJBwZABr2Xytf7l6k9JYgZSbtJZR1KECb7sR1ZVm8ZsROikmKhKZbQ+o
ndJBnyoeFf4TEMLPScHbjBvjfzEQ2N7j3sJJ9748E+bI/YFGm+vEZ3NMYZziU1Ls6dMovl1c2dys
ppbm3bN5H0ZMgyEneCD3g3q4Hcr4I/bAnz+zgZOsNd1nwWpgqlQYNk9TsxMfhUxOPH/wCvLHouZ1
MdoaB62Ggb/0tqCFWkPfEizMHKSlSwwI90TjjeMWHGb8S+CMNq46R9tAXFMKoDRiIegbJOJVRc16
minB/jy1inenZweLJPuE64drDecIZiVNfYhIb60fLhVNwwEX4/3/OBWbpQ9QCetT/2Q2Y7zxJiFP
7HlN697nm0w+aHFspBDnjG1+aV/4+FQwmlk2BJzvc1ZWNlL68LkiJ6RXW6CvIpuA4GCmAnIbjET1
vV1zEzWHpvT+Ks7VLGhuKTW+aDd67pzSpQkUhXUsr1GU4Jy75LbKMs48CDCvQYLe7xfU3LyT4ppk
djIgaNAsVTseJAks72k9HhfHrY4Lsszui0jaUol/95L5lwvsrFbMeellz0SfNX/IRuSwEgJQ5iFS
Tsb2W0CbAb+5iaPQc3Q1+kxFZCn1nJa2xMn5MvVwQWv5tmcds8y0YOeB6FQDCNRUy6R+GswLOkSm
/tVtSx4hIRysnDbhle65b5Y6LOa0U9yjdAmCGS+PUTr9RaHH9CkyN+bXmzdwHnJMH6raBnrHubVZ
QnXgEsjg+CgK6DT7YpXYCGVQ3RPItEWWHel5DoilnY0bmM1xmy8/Li0/LZ9Asn5hK0qXG6yswhUq
9Gnep2QgzXEncTfIBrBFvS+ktza6wnU/7bb6ONcgeVxrQMAM0b3eCkXuaku6V/xHkcmV7+RoHyiH
O3lGutvTck32/zZD6BjoSDtiFr5l2DwtWsl+jsBvIZ3axNsW4J3vZK1u+m3OU1KAM71wfYsZKY2y
oWy/e5UvAZg+fIeNQe8/JzGbT1H4b9SHoibHAfzqyhyyoZ3qNLuiT650evwWSXYqOzEEvtaccZUN
TMT2TR0LLwDlwTCs2JSoxCM/JWws2QFXL6xmfsHg4zmJnQ4iikqOWGOcZKrXuOLF0fs5afzCQfmJ
0kPU6uEeZkUllvpOntYdbPdhIAc1p89ex9hkzgLTNk/HIBxrSuERC51hUgxJL9hjEadK6EkNuY0B
ReeDRUVSKOHQl0HYpOSuK4hVIoXqod2pfZUOVedwlJDKfi64jFLt8n9oRBmr5fkNrLbnkAKoJMiK
NdZkceNSv6aWR3tnM8ymuEogljttccBXCu8Ezz1aXPjEsDPJXg19AqupCKMLHE9t2/If46K49kos
5hw/R0fJvUULH5DqQ8FWxAXMw4B03RSozvl6GOTohKfMusc3MwX9nUi5tgr2XDLiS9UkaxFXyCRh
GUvSc/uun7tQXN1o8r+FmIHTIA9zmGUGc2TDKqLfQl5Opm60TxDKKoxCen4T7UIGmb0zHPuaaJGh
8vO7bv3ixJxGxRhVssZYlyUXS9OiG9vs3Ly3UbM8/2Nchg77JLzRisx6nkQYEv3MihV/sfzhMU9a
bOkcd42Xa/rByhPSbVcSpd3dit2zEhJiFXiKEDIQ+PEri1JxERFtXLgI6TFAF+JcVJ4ccP+jTXs7
ASfbCn9EsEUnEGNXOnb3oDoeY74R5bDtyGRty9HkUDA28hBWDcuURc6fPEiEE6+pcqMNxM+LkirQ
QSbg+3J7wZCuIquV31L6DriEhgNYSJSHCxpkgRrbAXWitIV2Y7xKqUN8mFjayHKA5hD6antQp/Fi
d+q8a3kh5mtW+6t3DYKL/RRsh56iMZah9D/B+XqZUieEMYsA1ef9Y4k9o1NlJOozxoswlNdUbZvH
wBp/yf9HFN9F74/mgl3A5UqhdzbVAeEtuyAp+li2z0NuSawsUuuxdHv1bHaD9jbpUYH/3+3n7nVi
k8ATKMVnH0E3uRrUkwIBRVTdi7JyTiUGof99Uq/o26DcYrq9iN5M4sWN71gXTApYTZ08ZiLM4Yhi
wLFDqmYgjV+4NAgi5f526yf9SO2FRC2tuKtHlEXvu8k3lpbqSJa+qY88kiOkpHxhkSW4o9pP5wdB
dp3Pr82EgpL5tnNHdIiI+8uY1EberlwCOK48fjxhnQHdsgT5JF4IUu3R8QxwiYgVof6NNHoFXGTr
J7W5hJK5OLIC2WJjBWd7b4sProKx8ZRZT1eoSaJYwtqaRIy4tcXRyto/fBiw4sRqZSy+2tO6jG5X
dFLMks8XlEf6Irhf/IzI4JMLXxUK6WtGIjjs4R5e6QFeACSZ0l4toK5ax+GagrqypSaJsIKKB252
fj5gn8W2CxC8MB84ShFlY3RKNvq4/ruCkfxY9jnBTPh5c/F/YuUyzZ4T6mESuLFXra1RglZt4b0z
YRpN+JnXkjnt58ogzNyVu3AKW4QPUsABjC+rfedmg37zqymrVbHjFhTsJP9GhA7IOasm35C62W0S
yZ58f080kkc0kuOCUNfLo73koOLOClEb5mGfoIcXqRsDyj2r4+PdiS4yps35BLN5awxPOHIKgJyj
bp4Z1HjbuBYN49Rbubwu4U38cO9yPAvpfvXMlT3uxqtpjMuNi/+icmhddzmx9FI00es7qWuH0EC7
qOtC07m293ZqvA7W1+niRhEYu5bDpRVLMENZSQUxTEFdn+PlDp+lvppetlzvs95j8W+7VGtYaMHV
oYkNLRMjP8hDgO1SXlwbMxVG91Z0QJTwzmCFl40o0AaKj9zq3uNRM0WSQ8+HxW90aO1hsFzwR/Ms
R8E3pIMFDOw5GSM9EXugzzlmYvnxJP8ntH9Zbbe8KPPHUrPQO36wtUGx9b8LT0TOUCclHSHJcc6C
Z39IBvAoVI4Zj0IYKqVDX56gKn4BjDX+BUxWjGIL0y69LYtcEdqGnlp8iXa3JGBegvOUvw2470Uy
W5o4bs05z2bStE4JG+s/PKv2sQOXm4VTcCUXlRlnXUqDna7hE77rFM6G8jYbHhA9X3rm2d/eG+TV
SE1w/X3W+CsXJ+RJu4wGeWQTlj5Tfj5cWxlIpihimr/cSGzAO609cASR2+rZ1unIAfzNbuFKqUT/
M43J5/1iqVQSnozR2y0HPmwjarUBjq4jtBZRqyWfjYFZBkkuBlnamz7PbdQMIjjTGjoEcND+agIK
jEdUpbgka/HvmDMTMAgdf1I8iyrmjHVwKD+yY1QcFgdBz6AnHI5Lf4lHLL39n8M5thPeMoV2pJHA
o4qSXf/sPSqYopDRkAqoNetQcsKb0IyEj2+F/LHUKDThOQKGWYYZT1X1s5PVDl1an7NOL50a8bUZ
U/rOL+ce8mQQDYY2MuGPrh87IrNyDlst4folbPBFs63IyTurjeXBN2UYCXxdQQBBqAF5n3UHBb1a
VknFmIF4VR9vgpeqbd1rqjhE8fPrgLYztsZsaB6LnvlUxfckm/BqR/ThMiFTnI5GdNBACdTpyWZY
L9QupJGxZWFoQ0W2wo17GFF2IVBDOax+/os826/wGXjc4ZX4pSCkbf22mjwyNh0Zk+Dcsj4H+Uke
ml9GlxyCUFTuL3P9aJ0oySSPLQZKmPBmDhl3NSXtsWV1j1W9i7xp4EiHoTohiI6iPyHSoXJP4Bxc
Umk8fp2ulhjXWxMgMhzP3ebwMSecMvWBYpYZbcGUlIRIEL1MebgOdapmSx64WFUPm+PmOqs+gc2k
XTuYOb1v6+zyfDuL2dtHm7k0A3ZBJHYnReVRbqcMd17GHn5cLxeCdLyMT3hTerAVMGRwNTs86iuI
tZpynwlttItNAEED2sjp0UnkLc4YwlYV2B2cqAXq0jQKrIYpxXV8/sNWMgxrh0pDfn4kLMawgRv4
TcPbEGkjoyDWZwTsSKAonsAew2nAAChYstPaV5gdKG4p1MkMru8CPfcQJ/NHHcPp1NQ9Iv7gQhYg
70ypMmW+X+5v3Gx0pyeqMtqYTjQtyPerceh3wa66qNacG33g5mwlKuOlszrFjopIz3FZPp/VuUTO
rYG8xOmFVYNdNcmAsdMigtrukxmXkeTDu9A2sMhPrpFLOJSOD0VWndtARei+ZCi5eEKLxztHvme8
rVeqi2tgYVUc23bLHztT1KztCTj980EgL8sFH6fFY7gELmAfFPzgxFY8/esArKSclz78WICNpE+9
QkjOX43gXqGy6hKQMe80r4kNQ36C6DJZw+GBALX3YBCqsZFy4Co/J2s06bVOSDKbpyUR4N4TyJzP
zj5fSvEqrXHZTy44EYBWBcq8oHQBAFvLkn1fC5QC6qtET3a2qDJhUJoJzxLEMePfcxWwaqRyhBoy
i/OLqrn825ny4AH3y6RUle8JpCzQ6bEpfa7Pe5tpjJHFF+PTrLnZ9TeFdlO95XKFY3WAqA4sPALR
l+dZRk1oCuZXfDBkhIhS0EmuNUvrJAFqrZ07tJHwnvuTnV7gaFqxL0qP/4cfbsqLCUsKykDDnr2q
rTt8GvbPNJPJVPZF6AiEzDq/LTUeQN1RhsVt0T81NuKnTIa5hCvykr0o8roLUEiVZj2FPimG3VPn
R9txU37NyxGxWweU8XlStWiW3cl8O8BbTVsKviGiuuaiL4JsSP6Z7wHmGc4Y34x6tgYpWRR/yljf
BPJbVgFvbWhbYzZAy07rJQ0ST4iEfWIt0akse+9avZDiD96sJLCkCcBfyl/ExG0GcSepscT57DCd
2jxlZB8L3vr3AjJ/S/bR6UXBQO7VKmTVi/qCO1soRXwSSboJXp9UxRzqGG3ZiU/FnRbol6fsZg+y
VfSN5r2orFUNKqZQAILmW810RsnDSbdmyBhxfYhXrztjYxBBEXU1+IZI3d2GbIhdlrfYo6QMIXf0
bmba3uVh9v8vzvBhLWSBJY0WiUD2TUYpiw/RmCfVd+YI5oTcFqK2jTFzoaC7SsvAs00g9He3mywV
dIrckvFt2fOTdEQhlIpId2A5WJ8o4uBxkuLdMRFI9IRXCQME8xATTVAGzTSWA5ZTOg3Jpe14m42p
wrOw0abcItnElIn4Xdex0Bu14Et2MidjhCuHbIQgLMopLyRiWeMUQ/EDuGNTjQ8EwIaaz1cjKH88
4PTj3MmMGHGNGlo7qJXq9ugxy07jssf27k1AISp02GdjdDwfRqWP7nGLdJDTS/W/iPWq+3UTLM2S
ikPbiSigCArI26lu+he+WjtC4Pjjwt31IUJQDgNzJjUB/TzEmX1AjEjEWw4aDr6ZkdIhVhrJKK3J
/gXOo1h/FXWK9qlw4XUIScR89rj86zuPxesrKBeb4qhQSA7+D8WhzJ9sbe3I1q6DK5Z0fc6LZh3y
8Oc5HIQFzyiPXm2wg7v7kaY0qkDock1NwBbpqrKxAHjnXJT3s7notoeh4tslzdXAgV+OnNL1+4bf
VkvyY7d2hkWtMH8/jkz6vD0la4vr8CZatoZHEpxKlrjCjmgYJD+Rtek7blKIRWTHtlVmwDj5NXJh
sAq/AE9gSb3LTzecfE2kEd8WDNIeOiIXYdCm5jswnO0dSSZX5LqkACgQbXhFsjAHyvjf6eS3GczZ
Wnuzj8g7Bxa42EFu1X86fnJwTb/0xQIW7iLC4v85rTWetB5B2hBSxhh2cqe0MJeGJd6Ki7Q4aL5+
F6o5vSI7ZOIkKMPbomS5VFEDJhpfIA2BbvgQuoLGDQMBqtFepEY0yDMDA2vyq/o0D3OW466F5Pj9
tyAR7dADUOn7eAdXSqEg0PHsLemFPusTPCEcfK+/EK+pq1tCvw807IeFrUjLUoRdbdbFzbGjc+tL
bz/ACb1ySugbvFwDgU+/Dk2aP2BIqUa/vKP+cM6it0VO1hGEbIhwQyfEKZFvHSVNpR0atlljBWoI
esuBvtbamKrlX9a91RfmbfusraXgSAbnzyow9+VN7mbyH00sXwe2byPxZFzJbCVvpCPQWG9DO09q
F/oGv9LPRCRwcFdt6yXvRrWIJi9Hf1QkaVsNkBGAkNAcPgDteZdsTniqoPjWG1QINYcOYEj3Zh+c
E4OJstf4wQTeOJvUZ0RvnrXF/ZSPhP/kpIQp8KIdKSmtvCfK37801e0HP6je9EPmOKYNpSN7SDOK
5vMyqTh8hD/j6SxlFObS6Nr4UcuH4quRAhMi4ETj8383Cre0XeaVZ6lLLXvvS2ra7VwHe+LAomKJ
/np+uVqWAmIKcZCm+mLso4sJHR8J/pOSE7JkfgOLH5mG4tBE82hA05x21nVqWX8bO4vgpTtLjWuV
LV7RE5NLJyZxWhyNzk96VoODzF/iVOVgkvvM/To/lFB91BZvvYuzgKy5xmqZEL+BVvN3AiXLmllA
s+omQ0KhRTInhfD2VwbD/7+KtyZ2l/qoHAerTdmWkWBAxkKP8fO0XfHu7015HC7fuU8Rlf9sFsLe
gMVAlQQ/pjFNo7CO3i0yKoukhwjKPW5JpoBzMTYZlQoWcI4vLJw5cRHLfvW+HzygIjNP8Q3YuZ02
tmuMzA1kzUARtcWL93b/zE/i+lSA3t8lPaiM2UGZ2lDEI6mSc57OjD/aiZZbP9Vsg0K2/cL4paqP
LyDKntRVfJ4bvFfolX4s1aP6P3fjyDlpMYt05s/G7GOATZE5lO+cCX1Jxf8CFk42Js22NQrBXNSY
kY7kwd2pz1FXhaYMXLfOegurYlS1RY7odLsw9+F9K86a68HlRvQBR9K9C0uvuwlyzJXkEcwi349m
418Q6mRIPFRVpjZfEH0hASW671lUEcsr8eZ1fOZVUY+reqxCLYsVm6L2dL8RCrwsqqvShBdHI6J2
EYMPMSBWyw9TVocGQw1Lf252Mig7o7BveMjCZ/zwjln2VvzVsxPmXZikNxqfUHh+jPM2BLPrde7T
7V3caU4S8PhM0FtFmj2wTclKz5t/CHPtQnigyzNbbKjcoILkEWxyOSqtz7158u8MvH2bNywLgYb2
fIVMijipokfvqfas1E6wfhHbIs0u68dEnMWRQ1o1RWdwaZgzC+DWLhEvUh6Ek6wz4l6H+fh5xI9m
6gPmu0+WyoUyG5JnPNXHpZwl6Xjz76y2DSWdL57N47yXE1b+fgijjNePrZLuQNkhPQZIbQBmn81T
T0aPaLphQiJsqf06N5XL/bVccOF+uXUST2U+TIbH6puPwGDpqZvK+xJSVbjexlU9GvAjaHjkTe4M
yspASK3z6MrfacyVrieExM06PUS56vucN8xk6pRjuQFHGfBDbDwZu+ieROU2laWKTi7TCXJj/o0v
HTfHCiCjIgY7hYjSxkVg2hCWi2fZjc/o9wkfULanZxgEk82QuEQ0DyTfTk6bKt0X0BhalZCmGgzs
wt/rTAytD0LX5C0ycZ444+W95qfW+uLeauAXyX1xMCa6UCG7EAZVQiXsJ9tDxC1rWPoq/0lrjhV6
ZUezoIXr7lm/CJ2OcuiW4JP+H1ZbIQSj8oeXR8LNSHtMxVpsCt9IPrcJWR7Rjfe631J/QTG/AM5P
p94bvBmnp0gswFAO3e+3VTsnoA5c6Ov+Ws3vkPHrRZSPgI4C4r8jAdRfqR8ODQppBWxRdMZA4Tel
Mup1Wo8BXH2PZEJ73oZGWOaIDaWLjCjWIOcrk0w1i75VqLeW8EVstnwkX/p242XRGQ641AW5AoMm
3uUe+9OLvgZ9y6/HkjIoxGzxj6qLk3cxuZpcBjLMJWoo83hH+UH1Fi2kK/zhRmTij1wzQqoKg12x
K3re10CzIKsRUgsZ18SPXNg05BG/SeySa3sjv5BiUxCfV6FysnM2UsSvezze69X8aqzukyMotsQk
mbpOSsTa3vp/28XYeA/Alw4149+GUhP+3EHEqB2td3jIt/s0JfwxV1e7fJQTuF7tPqry1TFiWdVQ
9qxt5nJIH9TFvqNcdtVSOt9NfGmNjcvNqWymOtCFC+T10ICSKoDFazciycv2Y9DYEVDS8tajYF1z
cGOULdP7vq/vzX8cp+vRJxlJtEIYr4uap753acXYUSoRSSXjZz9YY7Hr6Q8Vp8SpZKkXNYAZwAzJ
W5zIep4eXCKJ+o6RLu31fzD5YIi8XMKF/Jaovntw2iWeZaHIZ9V2Dw+Fab/VZ0krnSP2r19WV4aJ
ivsHrpU5Fwpvd5KEANS1qkJmseEsbjCCvYyzb4i/JWUZzr6QwdyzGIPmWq0CKH0zqk7oIdZX3U4L
hKFgY/h8FJ6Gb38hKjj14EZcTOVGwebsxo6DHhmAK6SRNpHSU6bmPyyjj7v6HXlsC2sNLWTvLKHf
P0NoX7zbNC+ymyQqmou2krAnfww6/ByVqCe5XoTtZEBbjVnTXM0nnZCRMFHxps7GjoH4ZXpD5y/F
jM75xfpHKnvPHMUCOfAhjyhdqIPbaaKyVO110oJZ8koxFTX1KsGG6r3SdyKcuyuNwdxSryIOc2Lv
+GaMNNv04DzTNVT2fKdHSWlXGkUJeV9atIsPB7sdt7sz/Cxfui4xYlMzDxMcTMS8YQp5h9QmBCl5
YbgTOo/kM1vRmHFIA9FxZA1Hll5vWC7Mmx8VXKKHbMziXlfuADHEUvuTcPl5PIhv+q38ka+r4lCa
h6rw5xZmMn21zeGYHnUmZ42oQqtp/PzB9jbBM4QFM+oIy6sFIgm/0OkJe6/IoYyXvFPhGZP4cRjO
K6+yjF4pB90T3BzNxZYX1eg1dlvJUV6xgJzSRH1TgyY6CzOQle4NrK1Zh4CX18oAK5VHtB6uTquK
DoJocQNXL9AUMyrZ7LLdJs5ipl79oHBpNzTSWoTWIlURjBRgTRgpjqxhKf2pEJ4CkvntoQFad0VX
h8pcM1YAz6I8pG4P5sgWc+b0ByTufKnDWllojeclF4B6mxiv1aZwMxx+2AbXr43CjO0wmEzUA5y0
bL4SxRfFl0NgfNylHi1nY8SLaLb6q1nInIdwws239LPA9yln4l17Tuv6pYY41oIw2vtpvB1NXHYh
9p2lrgmJRACH9UR5HQWa1bBZb+fyBVl1cpWoT0r5ltHUMbe0Zke9jhNSpd7T+EzFquNI+77zpmze
EnYaiGPQ+XZieKZczl0zGTBePBE1Osae4WsgmXFeWUXqFp2e4jRNqwjGnVqLZmVuINHwyaJPTHib
BQc27QYCcyFVJzOb06XNAdBFXMpSa29IPL0remd6FTFe23r5n8PiWvlN7jFjR04VyP9DYIjq+Y8y
5fVxAhgf+qKO9/+hZy/fUVgb8GKVnJBBi7hSq5calkPpdiLKPoOhGfQ+kSYE2bRnDUmqs4tqdmJP
aVfbB7OISCDlkMvwr8ninTiWUYGqXUSy4wkyLBSW8U56lotwhr3jyPsiCMBYqD+hjiseTEGnSAhA
P1UFkIqq/KXCJ8r8HFEwTdjkZXf54pzZIjLwoaMENjyWqLg5NKQKFh0Hgtezt4M5tx/GORriFD9c
P5+gFzJLeZ6FpDRvKMDOMjnQGuKFCE3r3FW/dyPQheUWFB2ZxUvlEIm+wHFu7tYWfGnAvkk+X4zB
GlEwn3VCQWm1xV9RACD7Lx1tYEeCWsXYFuUNkOchfxNZF7wi8DWWBK031EBfM4kRSHfVR3mH+6Z+
FxgjD0okaMU45AsqMRdfXA8MhkYtQz2w4p2AIn3/yNthiwGelbLG/VhNasIONHTlcpGsxeysNCLJ
h2/qAw8ldoF1a+lmbeAFlsxc86TeGqCTXu+l62i7zNGkVbMOfTPJcRTT9bbb5vgIQNjAbMljHze4
trxnMNadC/6U6keLaUgNO5F6DaQbRY/bhC7S10JmNaOHFK7B/hXUErYX4x4Df3hsfXfP2HAiTxjs
gNqUmAY/W6IiY2ozDtnrTepsuYYTREe3vhE3wStuDCUYd+tvOZJWQWgS89GdrRS2INFgh1QCQXIw
rMkxDMbIt6bhgswn1Patr3sf55skmIAHABo83J8iwPRT5cm9948iYh9fRMS+M3812trufiQCsosM
re5a/6OEsp/uTNbFOyM0Y8wqj1urS0UqzHinr7ZFL+IRaa2iaepgR19ktS0PQjr0z7w2dUGjMaNA
BnuJRQQi4CAFIbxBNQrLn4L7FEr0GmFcF3zarw2rDrOi+E1XYQcD+HoFsQGwiDDRpLDY7hxucWXi
0n/9gODkpFeCiWEvG9Q5cIz+6bfsW4mjEVtq83SiSZDNqzHVUQLyRGN6f6saVvsR7I5xrWgOc9T/
77LFMLgJLLi5JJHqGQbI15QPvAax2iDCz53z9NcZf/GMJC/x+2bh05MIpdWe05evhs+g8QGCt3UN
zEdUD16Y8Q0IrKVzrwfCLDtjp9sEmw1A7/VeTdbF0mg6slTPqQt5v3Kim3FDiKLv9IGxp6mn33ww
aNehHYfZOpejCrBVHpEMM+AA50G35Hc4pRqfGdpsX0HtA+HS93VW/BIovGwZtz/kQRcDXz7mYpeI
AOmDBd7xm1lZSO8ieHLyNpxLez0XWqPagDN8p0ZtYogSEW17ccRcEDGt3foNCEqkcdkwZJVfQZ0r
OBSC5/GphEuJINogYRRTwejmkWfT+1wMQeCrM3jfVr+k2rAn+IdjxE1jX7O9MuZQnX7QMrnUvnwH
vDnx0lPeAJxL8yAxz4KVAYbzWWa43xTJWCxmfllIbxmrEWvLchDCNmp1b3pxqyhWfaWOrDVy6rKm
55d+yacwC4Wz9MppZyK4PGQNMVe4Z7WMsLuqKFb1P7bNRm5oyo4dx7gazOl8Wu24mfxHBdjVvfP/
r+NApg7LWOGDzdN3DPfRpdifDQM7wBzNbjCz5HP5xhztalEr49l0iu6AXzQ4fe4XM+fcdtz6Y2Rh
macOMz+UVYD4pY9npVgM1CJtZNUR83WnqUcekwt6ZlASGk2xejc2u1KMi+5N19OrjHn09XNfoUSZ
bgveuaAI+ffnGWxscV4Suy+BXPvsumtylCFHCQxoIbmvRTz/vYHUIVtUIeofj4kMykZOxZAJ3rRe
vbZWasWK3vrAuqaPX0zTVFvSDyW0847d56c+bpQQaqyjGvB74BTgCtjudLS9GRQEgfjZVxfKIBI5
/2KakLkRWGp79tt9d9L36bqXflAmHxEuLuGcujefRWxp8KxmDMnckcYihgt2JGfwOwDvkW5TSagq
zOB+nWCvHgR4Ay0nA05ypvJyn1WzYjrY9DmO4JPojPehzrI9mK2PK+4w5GZYOIRY9jwuKzeqrM/s
jC5KHVLxJFT+FZV/vZcUu9ircG3T/HOF3B89UeDxJNaqY9be6QuwC5oPwko74UCQ3IWqSppa93eD
S/DV5OdD6Daap7g3pD8+h2jxuUFfsoKevIN5DH1JgaYJGdsmd1PuLfzf9TShKRJPFOElkeV8k+Mc
NRslZbXwgfyZ+dA8IS1SMjryumrMFnCYwSwOuXg1skVxejhLYQHGWl+xx3/aASdxv61unN5FeFKV
GefPl5s6scxlm0DyNBAbpIdj2UYnDevR3uO1aWgLvXKl3EyjFfHkHUfvyMZhnFtL2ipkhy3wnRO7
9TdZFocX0Vz6RFnu7ZwsnC6TmXx1ihwFCRQm2v+0AcXGSB40WuGTY4ob2WbIqra+BWWmAJwK52kJ
u+VhDJhsspOTwEXVJ5koVOM4o63Opm+lHfShFdZEZ9ZN0M/bCNaNgyzFIoOO8z7qRu+JCq0aCAtM
AeS+C4qoHn/gDETZgXwyWdURta7S+pIttJbrRoapR32HCJkPtE0zEUqXxY0ct6X9SwEAg4d3ffyE
GHvUaLlb2IajVoK9QpVrFgcSDY/KTM1QZyOSwascJJ9etuzZmtHexELUiv6whhIiOBcFxakxTvre
6DqEimLCBh7zkFlaAWFkBrGmEwci8NhxeqGb1AiBEjJLEMLsyYHjCD86j4zlxbVL72am3vP7u4St
r6/YzrqvBBfZNs5VwhNDMfq0SbabrH1knAUt3CpTGYF+MXQ2I9OhcF74BMqZtiKc02CguHV0A0pQ
rzgabh8FPHG+IEpTGf7PKKgmRCGW5WC0hQacAHT3dRU3oFQ59xgRxDB4CAwgTvgONoerihvNPixg
4X2lRjzv4A090VYOFMo3d/MeHKfU9vRchomUyJ6sGSzJge8Gq+EhuXLE5xOtebP08xgq0k2jYy5A
hbjU1Ru8RKQKrkSvSmz/ohgkUHW1pE+lDGQhFSWVcIG+9iVvk2LktzzNDoaMqUXHJs5aIZjIk+V6
mmgzIy3D5nGJXQNhIf2FJLXyHu4LB/1xhB+Y0S1Hk5QYgKsFnUGmYX/jhgAiFu21430kDmLYULQV
VYCZQvrjA4yprwGz7kJdagEc5beZC9ii2DLBpmXzcFUBO/eANqfxIm5w87yoTlU++7jd/Bfk1Srm
SdmXphb0+4lt3tTwkqZwaM2QleGOzylDnJ6kP7ZZatXSrTjWVEhHvvES8jTOxS9EdkY5k6hN35ka
ql/hPuf+0lUVNVL2ca23j+BumTMK0mieDioeZQ7FmxOQyWTAILJoVR1UXzb+tumKfCklMGbGVxGg
CFR73z6fxX4HzyWnsuwkungBL7fo4KfISt/Y6NC2pHjr3vpNeHs67DY1zDFmBcO4T3VmY+xKaef6
cjUk/lJxnpeu14PH9xbykU2Ae8sfG1gfY+0bmftJZiSk3ByaaR6XZ8+nPeLKW2LZGcHlVZW5ltKP
n+9soHCuEJA8SYVmBp3mxgdyPEEXmxppOwoqZzJEakSn4bOjxQjJrfFU6s09XG7OeGyA5KJqyKCJ
CRXU2aKQEfXKeVtRc7OFwKGL+0tRKZhT74AK0FaBgUhkx05os5ZjgdZAuVghAWTSag6R+rnB0mCK
XUW4fL5UnTPS6tbKj1xfq7l9pmj+7k5LmkHdEIDejAwRtSC++CiWFVRcmOQ0T5Z0pyqZgXXKbA9b
yfQIYk+Zufd/jLI1raJkZw8iB0lbMeB8eB+V3fTlGKX6P3/0mC1sWWuc5fjONWuRO3JFnR5VipEa
D0GSYbESiURW9BZF0Vo0oIEh5BzgFuC8R/qRP4NHN6SEC9oloPCNGYLp+cSmd0JoJOxhjZ8KQm5p
m9MVkfud2L12RXGNMcAWwq/2I1uWhQUvs+S4Vs1LwrFBPCfihYOio3C9g/ygBrFTzHCF/Xs4qtDm
jZ8uRDDtof60+FIQU285zNtL1Yxg5E5sRmTSCkloYJPXucewfwtsPQf3R7TDPfnRgJ8ovJQqted3
ON7+g5+iufcrFmHCI5vQRj5rJMOleSnfxXBnfIEV2XIPxAUHQXUdKC8sMKgWFk0pcWVMx3IpV0Ka
ID6+I9mXcNIZVqA3Wi8WXtB48XkvgblkvZVlHMLTEAgguylqfDsp4DoWzvc+spN6xd62ZhBvc3cU
LzyYc+TC6NDGDKpcA5sVLxXI2+dqpiOJ6S+qJhDKfsNO9A2PB+JOf5D/BxMtMXcnuqOG8SuL/Nf/
NAULQu/Jkp1sfm1fGcAk42F8epk8+wbk37M6RamcqNokK6keUoF17wyp4bVZumxIv413p1Z/9pVy
0joX/7APz5FpWrrNi59ugRbRueLKEE6gDzxtGXOoNYbIl55HiiYm3OeZqcqCdhn+r9R0j4j4M4PX
Hw6QktV96pb/DS4GHGEK6W8+tWNWYNaj0VzwhF9SyFwfQbVEv1uaaY3Lwvs59NcmW8dXV3cAPG2z
0dLAFS7BR1F1DKZX8KS+XG/IE0BKJni3NEjjeHMRm9RmubGqCRxhRpo5rboxwiIwZv7HqOb0bBxw
yn1SLTbyu5ta9B0ogcNlP4kxZwRYg4uVZd73f/qPuiaBFAAdeK4T+WZiqcdn6XWHj7IAx2+0Ysb2
c2XYDhfTjI8/S0Y5QX4LjXF7DQBNK+h9T+q0tK/YGsbLWcfgAUFFfQXlnotuH+KS2Fnq3tZmQZbP
z1cvVJSdyBVJMMmm4mSP0dBPaiCGu6vSEhaVXgKd2ir8ohG5OE9RpHvksf8QuxrzP6VFRIPnTVwT
q5Brxue6ilVA+HsBo7TgonCPkJbIr7ILciYmAh6/27rTYIUhmxlBdlJr94hnR+7yhxbD/aKBtt3r
Nt+QKfXR5aVC3V1MvrhXfPbZEYcEBQ8G3aiofIUVQjjIky84K0pneYOR5gj08ycpdJ1kX2vOsdvw
0czgKLZS7ed45V3JUkG64BErJNg4RZw831gEERX08/QkOLggWbpc1vvyC5bqYeZJMxu6QjgWAjm5
2n9n7P+MWl31MCKA2nGfcCdtQRSjIagVQ4Uuv7E55HJFCQoElCle2InULa4LrP8LawirN7kp8JZH
n+eIO0OsmDlQEsXhmg7vAtKv7ssbNRKG6dZG4Sk1MB1nhRaf0Eay5trghYVkATUNvuv1Me4aUZUr
7zKn83b10UuC5wBVjavce457/eKhpfbNXOOldDHIT5aOZwn7uiOt/4RwvMStBvbWyAfZUDFpTx3T
Bnr2Z5Xt5l35tYNedJCGPWXUS/7sBchK/2YSJTEOzOWT2Yr4ozlYhT33gfW62BiI+vnZtSkHO56+
K6LKLdpKbbEDQXy1tAA+mHUTiX7WYfd0VynS0jBGCBhltzjdNAXXOxamljntZaXggjimG3ZaSDfJ
cdnx2sr5jbUctC7wRFGB3HX4kVFb5cT2yv8xu+sRGBvFTy6SxLfp4+iKy3mRUAQ5yiJKmYRbky1B
LrxSzHvEpCbH0ZrDXpaOkCNvk/4ySg2G+a00buqFIKXDhxfcz5ZmdculFkHi289Q0xtRizyJ9Ghz
CPJ7+OSrQnBQAZA1M3QVYsmio96IVt8uNx6de5l0hGXujIleJP4h1vpJ6h6rLc7Av5YX3VB5XYER
TK4CYeSqZo+DCNaksHSkDSpz/XvbxyZVoIR6BOPsACYlGwxvdhPWobUlrGZfPotPaXmr8Qt5T1sp
TYbxGSovpbcr2YQZJkcedL2x1TCHwXpme2wOPxHZe2g+u5Q66T/F6wJRmECChOxXCuq9vn3eIcZm
iV/Wi9vybAkTzFLgL21/YEMVRrn2bf3FwzvEp4Kx+l7fxhBOy9/efHcZ5/nqbIvoBzhb+Hx4c0dC
Cjq9btjlUdpu2FXhwNg9dsPYt0uPlrZ5yEdi56ekJuzHp8+h7wTJfiSVcUTf1ALEzkZ4ARhN+D7/
h72Ief4bxYalKXJEw00ujw034glAPKDsHmEuvRh6yJ2NfK8Hp39r6RrTK1Ns06+QV3efPQEbSppz
QcWJ3mArXhxDkZcIJ7UcvrtPl1d/CFCyOi24a40jhDZ//3d5H9Z4G7/dSH8X9uYeZdkurZyKTv+a
/GzxRc3u6FtBpCqFvZyowJ44kOvS3wiejbud2Cf21Ep9fOUSud29ud3otI3DZ0T9OzZBe7zvwxIn
SAU0aOx1lbbc9WIhwZSvelLFgjl7ZrNTXQMKwkAnUJEfCBL+tpiBt8PLiC2OIhsm55L1v8xIf+XZ
3O8BnymhQYMcLUBenpvs5pLzDaIv8r1WyToqkt4SveVzBg1ymjxkFBllc5RTqtCca91+Kkze/6Zu
gtqbIXn+M88ldtAr7ImTCYJqMKs0nw6PoACbUGXowrRqv9j/R/4NVebQL1lFpiZk4cUzTqRaKnjL
ZG0Ku66DRA+1CtIvhO4ubICzJBbugpD/ISeHhQ77p6+oYIXy/O/EuUp+G7Pjzh0ZV/QKu8ILZdQQ
eJdpil1SLAEZspVyJZ/GRiLwu/uPD4cR9zns8a7lZs0yyVmSWVgyl/5iRfXWOm9w7VLopm5/jU0i
OYepc7mhk5r4cGjVjOh333qF1UmzoL8H90Ma3IwgbYjOoYfd64vVz0tHLoUJaSAWmszUYHocZFHv
huj3hT1p33tsWbY3JZlYhhPddhntyPWWE3ux+M1X0kZifXCSfaiv+520kh0qtL3lB8Obnf48xOtO
jRqmLKx2Bt6/XQ/7TCaeoab1xLAwAE1TJ3S1Qc6ovfvr/inWsBXeuZZXVbdxitmRF11eAqqVKNIs
zoOy6mS37OM4wYf6+lnWl/MAjw/A9QvdiBhxChp6IYfARs5xwb5JlyxJhRbQx6ETOQAXYWap7rft
0e7gMAGwglfTNRFlgBg0bJJItYeg9IDETp2RUHpJUE4zBf9dfQF/0A7eaJEvOWDqx/9p9yW2RDpx
NV45eEOrZdHdisbAoLwSZs7ayWGYj+Vj+B609xLArioDhNxPCiG3FeprVU/YVh+iuL6fHQ1Y+WtD
og65m4bW4jfcq7S3TZdFnhNLyIqdpwXE3mSPWzDWAcX1hUgVWZOIJm2/+JpphzdaBotL37xXEtuO
cOaEB+zb+R9AADb/bE0q8p6sGZWjLlX5D2Cnd/HHwVOEkS00Uk0DZdf4QrkF6ZMcR/dgCnxYGNBE
MZFYhAKLuhvQx4uoVKI78EfWiB9iopfOTkhqZzfGyYpJj7/QlxJHxzWwpdRWqjlmM+ZTvF1EkFjd
/kfLBvmkski/zcmEkzXZX9dZPs8c5wiJdly9e+xPQ38+Kp6AK8/BibZzFNmcA+rEfQr8Ixml2qT4
bTEmQMbJRHzngEDYp8U8+YNN+DXtV7iOl4gTivMtYazYaZ35Qety7VT5wzP4bkrJWBk3svaF+Ysu
YBov8n2/sNh2U0IisRs3EYQaswddISg3oXGITPpHo+oD3C77qN5Ff9UgvwJNLICgQ/4S5S3cl2ZP
ENBfGwMo+jeYRkJWRryDCgmMzR5YIl62HNfrl3leYP07OFLv0cdzjuTPgseXcEuxR+xKzRUB7fyP
4RhBQEWUqzlldOZkvO/tW5JIxiLoftxLkgkQJddQysk4M3l7Em3q0oUlgd8n/jzOWtVk50JcV3Ij
eiLqSzd1FkvnijRC3Mkbp9GntaQTZq2nEQ77NE6OPFEGp8Yh8KAbDOpmPg26/okADfOpiu+MDIbE
TZfkyG+3EjLvw7d+04WqCW8cJzuiX9ACc8cU4ai0T1Pst/Lcpdn3Ne+Fc4wkpZ7tITIFTigiLSp7
zjEPekUBraz9vxsc5lJ96eTY2NK7YdsEvzMDv8DXK8Pa+dBHmGhn8F1qV9J1ERay5wEP1Fz1WlCj
bfEpUiiJr+DkvkEeGwurbZ+gbODXn3oPyEsfAMOpCajc5iV5GzEjXK+ANba8xUJLV8WaHQTkGNtl
tStRG1L36rq6GqrbCQNMc5VKGQUeTzOcZv+hPHtPNRZDpe9PRQItD/65PXUXieYlZSLltFUIq3Hd
r+hSCgWHmz7JspLuYiC1W9dY1rDjPD8Zjj4tiHegELyxQz9YrjcogL4k1+8h3x+FPaSva+Yh4Xa6
l0VC/zSkiDfeXxaRxOhVYyNmhO3RMQOaLLCL2fl204dyC8vbHJ9jYOqjsn8IoqgaEuX0M3BdrVqS
2ASBTvrnrjkr2oqvww8CV4/4U7uZph4B7jBoryLZ1kubrWhrCu92Hn0vblDi/YPrG6hL46y1rgvY
RgSauz+fnccZf6L8tBfQ3KjIY8+H/IiJGwSVset1j0WwV5po30da8v/XeRcX1D+BbVzGowE1K5CS
/XLrznSyhxuqmeFwxLqJGv57fdMy7XcsvgFaPzui/M7SvWVDNIcYFHOxQBE8CWP/1Drukgt2waEK
oe9d6Q72ZqKUmYxNuHLmFHUC7Z1RUzfBkfmoD079AzW9VVeuPbbRVbZdaxas1iU9k3oi98mN2ON3
/pRsPx7KEpeVYObzQrEqihs+o6/sFAZnNnAbD8oWdjMu005L+s5CofmeXnUaxqwjJeX+Ab+WCN7i
dzUQYouhat5hllmbKD9+uZwtrl20GF5QrKI6754AwWWR6j/uDL7TrrnA7JadnjiBZB8655/agpfL
2ceK92FzAe5kK2RztbBoTGyPaxdcXgxj5mY9wj6+GEuF3gfK1x3UhogGyKeJp+LH0VDBtr/mn3Ez
4o4OcNVo8cXmVE2Yhz+/8CPmDG02rMB1+bWkZ33ID6FOZy09tx9X1lHKx9w10arQdeL5gggff3M/
1fxg6yD5dYpxdJZOU+3yEruJrF71d0sf7rUOW9uLp58QjPjJVA9yiKE6VV8jaXggX+c8MnaoWw18
FmbDZDfe15dVD5fuSbW+RUIt+8UZCjGukDDSxnRv7j4PqAmHAXjxaB3cPtIuGnCq1WSInURa6cU/
k88ZXE4qH9gNEky8SmE2p80chh2/Rk+uIE1DBR7IZPgmc9xjsrU2vk/kBdMIFQX0hkiCcSveNJ1H
9bxslzcxNKkpXWLmY9331KJfENL2VaHg10TS1BZRUaKilIsWVsl8RuTRKEJdmXsYoBAC7aeH5d//
E/eianbmxJtOKbhj1c0BoYPGI0Gs5zvxCA2V1KD4puEYOAz53tYp2Q8q3aNy0byzjAjkUdfutrrR
1cKN0FRUqKdb0VhYV4rm4Nu6z1Ne6mB3k1bBwyKrcNQ5UXHnyOnMmnBem3cYH/dhGBARurL024Rl
CGmdZHkimrLffDzlWbj+YN/CLBvG0r0Y1Z5xwXUCY8HQ7s8PmEuTJxY+DPczm6gEIfFL7GSygMCT
5AXg2VBh7djtFlHYj/0P+0YeDsA2i18mqlRTLnJzMviujcnz6jgzectHnn1Avtr2wlGv0N9w7IBj
BjRdCz/YcAaeQ4xxqpa5nzQ5kuMVZK9XC40/37ScztFgpXBYgCZCsTlyw8TG/U8KM15tf8yzsmn8
a0b/T4WiudGMJmPzYyLzG6qucplJzOM6kreIJSidNlFM4RQBK5BUkA8SUhhqasvTor3c5nVK4trL
ctG/WinVNGBOWoZU97Hx7w6k1TLA+TOk5FtFbHmQPHcg2yAXk8rIl7IDk1Lpf4Zy/8q6SE1KpxaZ
g6ZapKIVDdANWuP7r6k1mxvTHSNB/iz7+oxDtigvxL8nBOh6BnNK7/fHaP4gwEID6CAMzZkHY8jp
Z84solGkzvLGP8iYzG+9oxYHbQ6u5Ak3PSGCdPXWe2yCZTd4nT6mk10km3AePNmKtsr1dYc+Pj9Z
igTBthMYTvHivhk/otQ97ZRe4cuQ2sj18K5B/fGLM1QX0VXXuy8M1ErqFox5GwbUVm8+w96O1314
UjlkgmzBdAiqEEp8m3h4r/6KQ2PG7gFVbZj5xzZl9t/7q+ksJhkmnQ1kNZyg4yHw4fhGewIlv38n
Adu7MUBVrNc43DLgUOnjIYCy9Q7L5PO0WoFIS9OLstVrdWFBTbnuIB/zN6lwweX/QSgzvR3n4amf
X2qaeKQmQZ+BJLqSZGV6zvPVqYodJULseBn6VmC+MQS6ZGaHNSnUoOrDI/sMHPyehBRRr+FbKMVR
0B/xC0MmQgCsDr4NNU85leihqPvdJaj0+EUPxFG6T1nDhPYxrd95n2OkYgIE5Q+znEQjmqAoc5bN
tOaaj2bsl3SdyFMB62sXF1JB+oG4VV/dz5A3VtQWU5qZnbgwIcEkLHIYvv+5rDUtZ63f1xVSGsyY
fW3KCvrN9IeQvjYJUwHpuQevj7XHvc6Jg4UWo/Fy0n2WD6zU2DVCZu9uSywi6yRgVPGCpAtIpOKT
fk8hv2tuow7U2iduyFg0Xzpxnr3yLsRS4FN82jbHeB6XNuPC9rVlxvt4+u4oUY8i1ZirMZV2Hkf6
mYHuBHCn9eC82ZOrIyH2ckvES6teDR6okEMMLlmGbPL+VCjAd5HWNemzZXDs27OVwUgoWbZ9ixk1
BuGSxpVBH/GBht0VuGf6rKcpuZhr6nzoxfv9kK/xaAzSAG+DIEMV5wgX/r0kwvAtznlkl6tp7B0j
Efyc7Je4VvHohZloosWI/u+Nt1EL8ZmS2pSUvpvBF7j3nystsuMgbh4VnHo4rBj9bj7pi8bkUfiC
sRzgDZ63IrQZw+/QbmzEMTbo9k5W5iVGTR0BZDlhrONzJ9Qo259ywf7N4CEBQNaZndzAbqlh8XR+
ggrU8VbVRQ0zUNKPemqvLXwEsVkxHwtAFtFcBLE4bmJlN/a/q8JPy/zE657jBWLDl8YE7JdYIPnT
NZLgELJgBzBi+Z453vz6tsM/DFiI/ZvyxMSWahsS7HnMnCizKFqpf/ntmtx5MPc4pK5+aZZwJ8Ym
djDAFu317EKNcsMtAy3NbX4jZyqOzUHFp9Vxc2WcBTRWbsCreuUvpHFNQwt+uuJC41+Jmp2MlS+3
gYiOIQJkWWhbITys14WNNORQ648jYANN9ob0b8vj5NnJ0/HDLXzcUYjr+t99B+nbFbZYkzGUVKZD
UuExJf1mIwJ7Qj+QFYozQeHo4AiF1SN6VVOiyAl0m/i1Iyuz3EVNM1pSL5u7nY1b0ax/lsJZQnNV
yObAFJaIj3OnJst4GYr9aLx39qFLTvba601Sgo0h2jIBdGaqmJvlxDxJsjg8Qj0YjBZJXWhXPFT1
GuytfKdF5z5RfsqJ/C/ks/PwM94XeNH8+XShYHM86n78WYKtncACQp29tv1cdZeDWi/0NJ1Lwc6V
KyKaDOaMNlAjdT2je/yrgWI8e7sI0a/g/4VaGTMd8NTMpAColBcht1jEkA3D/2g+lj7OLFcV7jC1
6gCcBzNxzOWc4blvaydyxTsXFsoOcRQHMXk8QNwJAE1CpirAMWXyqkcrBxm4a9OQNkUgPHXOPmYH
e/Z1p8gmn4CR+nGds7AOZh5eXpAyirrtnnfgXNRxh3+8LuGROxPRejDZsfnjMw41fCUgRwL4WUg9
AHUWeBam5ppn6Vl2Zi3bGBZe7N9yIdoX9frCZWdrutAQR1fJqfu+BYMAt7cCw23a9fQbmpzvuEtB
dOiZzoA8it/LLnXJ+QxaT2FzWPPq9ZEtz5X67jrgkeiDTyYGFMLAxlyPI+EIhTD2SB4snZbp17nx
xJcrsgJkU4+jGJZKdhm2SeR5ip8gBxB5FkPBvpuNT5Q1jbFm7u2OoukuSA9Nf2UO0bfYUju6M2nM
glE/3A2yJDU6sbHq/Rpr1WGhVazC/eN9Ad+uxuSjZmaN8Yk9lXJzs1j/zZvNyCVLXnAaASrhg68g
teD+hUfXEmfV4WDIq+0imZKqro9/a9aFUhjjKJm2xx8LULf7CCieyPysGd87svkLW5FJMG8cgU6z
wQ6kegUDgSXaXQuJ8QfTPzHcngk1j9tNzkm9pf3b5N69gbE8xj+3fPBBkH9FEZmCrmBgoADBFsTe
kLNh3b5qfLaBufZPlEBvxbRLZ154MySJBOToUWhUqJTZzEyhuxERjejmSgO4sF2u4Ju/cZtEG/J3
E60LW5MRpn34oaZqj85EcxHLF3wx74O7+olYUXaSsACxowQ8/FZ+WqTBZNYG5yjTiNYWvwsxIYWK
xM3S3BSVHB/nrxj8pCdG5VaQ9d0wNqEZmflDRT28mcRICrqnrAimZ2y48lSmXJdoca6TVVGOzES9
EutR+inoUum/Cgeq9ZizYhQHMfsg15TfPDLsxMJtd2+0p0NzACfTwLl7oKCDpQT2ZrFEG07RxK49
mTEsu+/UYmC7lrKKUrkE2yPLA2D4I8k8tVpVem3Mq39WIXBCyXVO1mA/sHJOnDUdm6L4GEEOahXS
qc4Q1Bkjd+D8KXS2v4tfpLtcsd2ndiK3dByfK+7L1zCPgs+uuECWXIlO7/fJK2LpZe1+3lekQv2y
q2Qee/Jvci+zVysOEm6x8Mi9zoz3DBkjkoW9rTFWpJsPh0CJSEdzLeUEBAeZph/0NFIX46y6JRKQ
5RIr+Zpnn2qcMv3E8ScGjYpqmk32DFDLoBDLyqOn+SfDOtzjy3SKvISTVXmCG26gsod/u6Bpng1v
l/2LZqeXpMpZoR4KEu+QxU4T8CtQB5osMca17/ICelJaPBW3xSSL9ND+4g7IR7GRl+EFDHXZm7Wc
6jLOL/YQPZ6mTB3NNGUIgOa03/nBpLldvmAHjkSepnEAy+CWcDcCFwoJzh0i1kE2p2W7G9kbvaTM
2BcnHDfe7HoYSf+o9AKxCcLPg7vXLTIGPk5SM5o34c/qPnQnt7ZtHygH8zswVN2wnGL20XcCNZgX
waLJiQsYGasn99MGmwQrUAdiJ8mBPuUwsgDvAWrkunnrvw9VrXKOnBZf5FFEbn/uZ687caNYQKYJ
Fu6GHUikQD7ki/aEFVmiK/mZaBbHHXS5NV0M/vhxgQ4rm57Jv/T3vRLm1LaFd0bx/I3h/ydKwStu
rnbQ1W2FBV+SD3lFuEfAe+YcFvdNANw53FfH2lz4cxN4fR7iIV6zeiV9RYM4DEfvM2+P+gmgUXkg
r0cWlxK9RcZMW9bSc0HL00zs4rozSUULjBRqllyc8jnIE6fkmD+R0rYHs04+u2SxsL1ekEwcrk6z
/HlKm3+77PsqRvSJ+dKK2cP+KBO5w2Z9qiS9gNFTdJIqvYcKQd7rm+8d9LXI2fdgVUW2BIjvjlwt
l7YD8hAIoJOtp5fbicUo/phZSNobxQIw+DPC+Ctmuay0uzDj2WN9A8gVylxNWHMf4TrNmzpBm1vG
393pJrp6ss1sc9sz2Utbw177nY1QTEY4t6Q+8tmAORjNJQrD1kdtV7DjxDjO2242k725YlYdLwdP
H2zPqKCxRYJguroyPFVRjSK7dKWvP+aKCDFHpn+F5PXq1rvB8zc3l2IGpyj7VMNrwS/5N0uMjBYE
G73d8cHzo9ZJl+IRCDYJgyiw/Dt5/P0S32BjQ6Xi813D+GJrvxe3pGcfVn85Vs93yjN2Kdl46c8p
nvnF0S7J3EnK4ssmaz1SfDVtwDgRMe0dcjcSLpI7S2S1rPeBjMZT9MJPh8c2dwBHNSyjytHuwZns
OP12vG4Eb4vgdMyIeWvc0yUfaWKdxuE86uMJ+t19F4KXZW2HKi2/5VJHEPNi7V9spdkq3KZOENK3
H5+v0NciEkf+646vcSrn4DDybNxE5iExTBCQD8BfhaBUhq+2sgBiW9Dd76fPfwz+xDbpVMZhA2Ag
bGVEG6UUoNBIlSvtk0LnZZkjdUaqfiKBrmsHG8wIz5fgJI/wk8M7dAeM3JnmeK2rFrDsAIVR+uEv
TB6od0ExJ3pGyVBkWs3eMqGBhvRp8xV/gwj8zA4+ttbayewBXIIxzGZQySIW2dBRHb4+9vtNPZhT
XQRlfLpAVd6w2uAmfYsfk2SPqlXph1ySisV2/zDHPsWxSbCnrll3KELqM2GT7fDpOQNePP1DyZvE
HGwn2Mh2OnqTrVdoeZwBSiJuBz14A3z+3ZBhdXExc9d5Cis4gi6sYfpnvKFiyBrmKhrocPkD2cgo
6WIPsK4jjd9QRoWnxvCZM+cpiqfoTtYaF1K/NT5J6X7pfk0gdsEhtYJEV05T39TPkNrq6p2qvY9S
JI7oBrK0JLpWI5F6VWYmb3BSHX7HnR7sFDjxpNun9paD5ScZZvRMugivT2PaFeUdSZ9GJa7R1zpf
b/4LDHlMsXvzNRtr4D34C5VBKNUnIhcqcLaxap/1C7AyAUCR/DjlWOHFIBVVmgq6D7VgumorAFJN
sdj71jVS4d3rKBn3Rb7LTzD7jFh/p4a+E9s9pNuK875hjrmSjaG0egZYyZGOYADzPxZORk3ftVjH
klrHR80J2Tx7Sazk/ibTaVpF7PX4r7gMvRs+SK2HrZIfkz3xcOajcFc69VPd5/SdzPqh/gQyDMb8
nN8QkMKVJ8jIqpBV6yt62bxBQTTJi4mTV3jsOMH1rhOyHzztXRncCsm47I2cGHsDm37d9vfnc0oE
TyxSFjX03p59aWBHHiUghqHVERwyrGMza2DLb0Bb5lPOQnScjFcJRZ8uOPjdDpE647wZSKzbaR0o
+4F51BANP4fxKaKK80AlWpaiHvgkrujh9evs+5kr9PTLu/3kj4UW7VaLuWylUPAKJee9ujSVfS2E
aXzygXi6CgT+IJpnQ5MoybFtNXztrF6BSz4MJMJvM9xgmjJ60MaB1S0ZO/HAnzBddgSOFdtPodP9
0hxJGgZAdD4W79iOj1AAZ4g+H3h28Apy1SrEwlTabQHY3TfQsMxp+FQ0JYkMsfmVeCq0tKX8J7fV
fvYtAQjcHx23F+oFZPh3z4Oe+CZPsJqnFmsmofyiXxCdMN+Y/i787L9AjHFA4CSYpdcMiRLixUb6
m57IoxMjMwat6dM7jie+FabReYW0xzVrkW1vBCkySacVIb8k5PJZvepIVq8LKzOeMCrkrfbhNxEl
GCXrq+kEEnpIAYxpEi6PVrA1djsqp1BTi1Igwxg3P4MZIpsLVBlZA8BhK3QnKCbu8rGLMJOLSepW
yb59pC5F54leueGSZgrIx19fdVJeJ01PUcAyiUWKlYdF2eWalNacvdEgsG5T+o7jAQKhIdCSCQI+
VgJVyt0PukJdssWL96WDomhzWkXPXIdtWgblfc4srzIVhosvYlHI0CBhWDYSYZXe3kvZggREuNV0
1Y71N0EM0PNIFjvvMmg7YMbRBJDDhWes6TxhqSpiSGr7jmivYYEPP+gMNpDT+borjTpHKszClIg2
h4Gfu64847K+gnJm7rPLDo83zNB4p/C+SIosoq4rLzCNkqxqguWTVerWzvgX8sgpi8eOzdPBS1/o
r2QKp/ddSzzh6MVd9LnfuJDzHMqfV7+xB1T8n5watACuzGK0hb3VUZAYpeF8HD5KFfweaV2ImcQa
w94RO+2COX4ilLUT9IGlrhEn/QwhlhM6AuRiek4KfWZYUzK3XPr2G4bejINhEqNKfiTOmNXBmxZ0
P7V+H6pT5D/zUbB0scmEUsKXdkZP0onS5ZDcRUK53vMb4OqTXSmRhwAidtAEp/tMUhpaLqTV6JEH
mwnEddU1gFAvQqaQ1JJvOO6DCPGT/mN6wIq8HX4t7eTK6RzmCCb1QxTAMCU4/Fxen/wTCJtfZbyw
YzwBD/ylxO63iC+PBx/0bC+5+DcmOe5LxNo/wwwFwXjP5YWK9no6EPTbVHrrn972ptgUbraIP5PX
DjXRwxpYkwNGiM8CAzLpU0b/gE6OUNjhQB+EmVFaulZqskq3oTGDRBEBYSUkDPd+QoWILOBpJjL/
0POzUYToZa5L4MrEkZBltyk5yWHmqhxIxOGorPxZG1CACNNZdI2dmQRv/wbdb5N+i2e7QosIFusZ
vdeIWdbDcRg1I8M5e//ozSzKSAxjCpGLcsADxllIaaeXaX6G7XGzXmUt/aoNk4BiyiA5uKgzxBMB
wmvPatLwLA7sm0K3rH6hz2Z8SwUv/XjxhF19WdAcmpMvmsz6gn5O0m+iSDWbeTJEUDfH8vAlk220
2skwywnBMqzexInS8O61y4kE2jP3tuNS/W4Y5CUFwRdDmw8SsBwkN0GN5yYxc7wTeAiu1qsQQJAG
78evyHuv6Dou1lh82xImsayvXOFUSEcCgHnOmy68sn1SZ8eYineCbte8HG4oTUBVfEOY8ekOgF+T
6iN8xK52mRWK0363bKmqzvGVm0g2xjTguEYMEx5VkouGlW9Icv8tQ1t0wmyuhlBSakVRkczJwOYM
c/6Ks4g3d54GNDGe5dHei6MkMirRp4ciKZ1xWNSnCnnoOPpmvRAWxkNrgD2/zKAweWFNDmY08oUl
CnekpN1aAyQIPLNx8HPvLr8Iejf/33vSa4i5058Vc51BqQEOcVXu96HxuBVVibFJU1d3nITXQRUM
wAWpFqKTVTQt+Ifs1bQdQ+NhvaEeckkK36klTc9DAZVBYMJ43PXOfbYKtrRroB40w/cX4jF7c0FR
6QDnboEPftQUnjfbnt5E16Rj1Sga9hnxQyXdqkin9JUnLZ8RcEwmuX58qyM0STAkq/5LAAFyc3uN
jxhVKWjyTA8KJXGDdkZYXZW00j3k0/x91kdPmkjxGssy1cX+mAnoR4gtAu9keoXAORgszwuPth5t
u+o3hNBDlSKtjPgqRrzSiNP8XAERIc7UR6Ah6VSSdNbQVpUJ2hs6PYu2/16KV/37Si/qI4pdCpKR
wXD+MI5hidXRjKccij2oBcLCJj7bvnG7tx/vIJWDbTHr5h+1P6dqPehI0svQ/+lrUxMYMicsog8O
/HEFHYzlOncTfbvwIpEgBWad2TrxUY/eDfkiaUqzJxEvIMcTgtlHxhKyJ1umMMyR2VM7Kcsqebod
8D+YkJiI9NSMfMX3Xal7Zx5ufjunAXVbX+ypUaz9NVcLJUN8RvTQhLx550twN4/R+uhn5cnfXU5C
qJvgGTEwQ+Gq32jJB0D1pZ18HJGHXXlrJUj+CNKWxAotOPm4zx0twYZ2mtE9GLTQymAIJWTVi6Xc
MU4JtjZZWJi+1GAoLI4UEWfrmtE1m1GIvFYWN9dLxhO5tAjQwV1TxFJvTGT5y3gjClAYB8xF3oFP
mk8lVuTvdjoxlSAJJT+9dFZkSaHIwGkDHIXWqZTIOfX3TSnMMY1yQOv7CDDkEt/SiMe5SzCNLkUy
/Z1ak2x9TLRXrxPdOUuMiz1KhCC2EfwZC67FlQOUg6/KuidZJODnSicr6GMJaH6822KmpE4z5kum
FhB3mlMpH90CnFu+E/5CCsPrdIZ85VbdsQTek7utup72G/CP6EQrUygh/2rwcDFAoe8mjHrvxEWF
Y4lQiHmB7leeDvfQgRhmqH2spfQ9xxisj17DKBUbhtiIx2B0IgXHL/yF97U3AfSWxwqS0gRq5V8b
G5ESW3I8uE3x8HvQdwzQBQqMpg2c+fqjXEtJJyhi/wXmg8bHdoUwJDiPqjUO5tvQqjMOMiDiirmg
uyQRKbDkjxTthtPsU8EwJPnd5nY8Uls95la/gtBd2bNcDR168NhLbXbrj/RZD+cYuOBAsGiuGf3M
KZHaAyaGWrfyqJ2yVyTWubeGXKHVovUY+PWSb7RZYqpFvuV03II8TEzH6WuhwjlLrpHO8jCuEdAQ
kS9OSIWQJ91vYiFkgtypgr9XPpNwSgqOuN8YVENgVKEXKHXEGiqA6JDdMSgZ1zY9lFkWiBGWJbDg
Tutb/GkW8wcSS5QBiT8U/3vEeVVSUrvmGFqkS0Vrl+ubakAB0I4vdAuFVC/YyC0XXVl6Q5kDJNIA
ogfeU/ItaXTzCttdmiHiSBavzKDYMDNNkHlTrRrrQDq0tPKXWwDsAlgibFdYa8S2WgZz+unLMRgR
AnvmnipaHrdY61oipxUEt8QUg4WD4QE9zgqBlCsNHmMa5caLYrFUfs25wQ15pCG5C3kxBfzlAcly
yQ4w0dpQjJBqC3zlVJ4QNWTI3OH0PbkUUFrm1fRNDzI222YZlg4iFlRJh6NJSYPiSaxFRColEsfv
66aXL3aChHREONX25HnjT3Ca/qRvmQSKLNZFuZZchdLLSElfSs4fBPeqb72s/AWC+MEdFHGxwfks
tg+CbOWPAHAcdbIbry5vXakyMVLXYGu8GuvvwuGZRSxGsJOgBAh9TSUB589xM0HG83IBMIIeyUIu
hkQt5Exg9/vc1gdigX2T+4DYEFbP4Y1/f/FNt7hsuapFmwowI4JSsep6Uei/XIClp1QsnKrJJoBE
KT13ioam3RccE890W0ADJWzqKWVQqyeCiSmKWQOPuJPb6mZ+AAfAqdHaiaJcZEb5uAfk/2ld6kNz
Z/MRgU22TZxPTyqeX3T7xG2JAKJ7lcfosFktLQmcNBgQQadIWtBEIq1Qvy4Gws1hlUA63fJW5luS
t70EiwAJPSg2O2Y7VqyeV8B5SuNm9tmyAnhqtPzWO6vEvTcU08yvoEfrLKL1L2qR3erVXtvDq7um
lqePCy3x+zAF2hvLGANA7N/KSMuqzC3umUuU+SVIAPc+IU7nhSPowFCS7hF26FIDGhNOhuXLHZzr
Wrj3nz0q6gR+auKTjQo4E6DHkYl0/d2po96a+WyN4xInzIO2SXIU2877vkwLgndYXd2mydFy/0cC
03OzPg0nyFh460DxUJIv4bI+z0ng7m+qoW4/KsbEpvCM34cpVE3kZWJ654T58FbK1+CdlhWdNakq
LTtrT5Dbj9miWOTRuskPiL65VUA2ObGU+wqH6mfLOwFRPJpW6Gj9oR3ZqvmPOlMrHA7dAnyNL8HZ
C9yYaKg+eg4ejKv9J6T4F/VuyC33DCh5E9GVnL4B8bMtvWco6oSaDdRNQ6IDBtXLF+QvemxGRPPp
eg9BvDD6HuzvO8qPvjU/dgPy6rQngTCQfLHq5zTxZgtyJto9xflc+5oD16XoJgBRAEdAn4UdFFYT
np1PyuFG/7srm0k39VmYe3Y+FUukImlWRLgBU4RaJDpoi0Dsm2CiQiM8kli2J6cwojtCvumgaKnu
IpI2Ms6GwObF6XcXxEERlduDxe3ruRpxBRifgnNL7DTMLB4aY+p0cIPsZhQketYbGIMIaAd2l6wS
Zk5LBWIsVkhY+uhXNvKm2Jz56eBQ2K53yOxJ4Urd6g3kN0oBqC9C0Q0DoLEwMnl8LsbxpouMeMXV
gv6kjM7vjy225tb/uUrigJsekgiaLkNgyOSANSG8qQQyx4xyxjg6PFFyM/SPMT77IQ9ieRd7jVc1
W3B9fb+NJ0KfVGXcLkeyoxV5aFxthc6PaR35lxfFxqk07J5sG+SN5L/lfNiMTKXELPFiDVKAtgDK
X2RysuT0/q94uE+qXZOMWnQPiSruY/22bcLLfe80xWTAYuM3v/O+/pfby190CcEOVzEKiIk6aGwM
bkSo3jNqoZQegzEgegAawPpK15lxB5qg3ER0dAsWXkFrLpKQ4FHh4GaBkkJeFA+yuONw35W8yz6v
nBvsXBR7Kfvilgn3Kw7LeD8S3tF2+vfSfIxgIwC2YCfdK2yPTE7rqacsDEmDiXvy526SOw+cbGYJ
84vAzgLa9bib8eBusfnIvaHw4wfYkaWctYwyxgypB2Zy5Eu0HuF7a+kq47LUIq6m6I03rPl2thsZ
U5vIXvyzWUlwA6ZeXXwFr0mIcbWL8tlTKlJY0ryJwEOAY0/cLgy5/OjYqIroBobKDTDoj7OCRe/Z
ZOusJPwlYBS7zrylkM675U8+td82bAPXvjg6CtQfJR29aw8IKw2JhdWskbAHnXPHRUqFyyU2jqaH
zDlkT1ARCA/V9sJgvP/mF+Q0cDcgZfsEIPHbXGd0+Fj+yy9jpzd6hspib71FpA64bpmBYZMU6EEp
Ius80ToQXYAhLHavlpV7RrQTbJ7IEVyP+szoOBePLM8gB2NVFdDTY+Q9XMMnjrRiPQr+D4e07nAK
hTuR3mxcS6V34pahbusomw154qz6u0t4Ozt2S6IgufMYbpD9izpxuSHBpFtfhDPuvoJCytT8vztY
s8Ep2vAX/BrZj20f6sdNPjqasqPAjU29NFJi0GEaglH8DDzofvjYukFsymMe4EDbvlsSDzTQBVGk
XLdimY0BMqcgfx6Oo4z4hEEW71jbrmIEy7D/pjDO0Bz/9PL3OruAe9gGBGI4d6y5Fnx/EBbB+8hF
MFHhRZwxPDnSNTUjPYsqoHIoaJ2I8uAIxqAfqAWEmnBydyb09xdQZIRipV8UVMIDEb8jDh4iZAfb
a5AuKcsz1NTF1VK0FtNl6EGJI8oE9kgY3i5cMolUv9I3kp0ZegRcm3q1D7c1VSNNPxOEfd9U0ieP
ioUuF1anEOnXQfD1W6h1BoRIQCIdvxIxH3ewdISOHExv2QFeswo++sf0NAsXg0qB0u3g7ZP/mmbE
Gph/nTocuuR30fKvLKZyn3N7RMOrERd16QOx5JZSRGLjWphPCxjpElWbK4ZTnr/wP4wj240qs3A+
O2R8tWEiEP+1o/nPhHtTBDM6HKS8rugYtAN2nxYz4O7Q4hXqYVHXlGyhGnBdcqaSJo3RizN6cT8v
8c/kzTDP+Ktt0ZlPNGvNgR2HtLszlYnnKb+dVPGVAHv5Pr7FTLHcGgmkd0uIwqazPvSEIuc7PmXW
arOY1AzkDZ/O/RVh21tlW/pHGHkPyH8A8MltQtzhIXLCw4vwakRILcL0w03G20Lrw7YpYcGw8EdV
sZ/fvgs86kobXUNXcrNi5OsmOjVDlaI+OJ9mcKIcee1CZjR6XXck+0sul5X8tNGr7DMVIk9SyNKu
PCpplD22kG8Srs6CpnkfG1Qp2SdCNO4p9t35rLOdqMIThN9lpMmncnTd4s50hHkBwG8stVfd2FWN
A/NWyiR1BjP5iVjhwqkHD6qHqO77x6DV8nOBsprxxwNpeVSO3byN40/fr4bBNzYMAK81LqxToGkn
9R9Fb0lPpYQj0argw6VwYUTiSyUBoxCN9f6FBw6Zctwlo2mgkoYqp9rsv7aV6hnVAy+dNNYpYrZj
dq6UR20NPM03jWd7OxVMQCSCVPqOpujfxn/hr1DCWtvicOCOmSSLHec4+g+Wpef61x7XWKsSSaxc
TeAQOCausAS+6nFaiRF1SO6gVIBEDKC2WDMJ5xMd/Ogv7FMTzg8WzA9AOAxKUybGc1OcEDshiojg
NS0CPHlox/x6Q7QDYTNKfe/mtqreWHk9XQlZ9/oZCdKRTui0n1DBJbaFyFGd5GSo98eFJoOZcCWP
PDPk/YL/nrIU7oPjSKsZnzZnGBX/FSzowzjrUIt9Fqrg6lt3U7+yW/BKMmgDJtE6RBb1UkTVK6D0
IUHuloGxxLIP1QciGll3fCGTFjuecxkpDO3gqdARUWZtURszk7W7MqDuY+RD2TttXhfOY+nyvQDF
8a/MlIZA3SY/+qP46z9ChKtLyfWO4PbSkYX8p+RvtmDdw69fMKCAiXStrokMPvADvPhH4YnJu34A
+V/p31N1o5T8jyNJkuhAqvhKswP+2pFpoxliRHlPO4YHHa5sSpLb4k8uaxipgWReJf8UxGDOnUw9
3aK2VHH97gh6xUrGrq7OCZRy9mmc+NawnR0jRJ4mkoznvu7S7j6/BH3RHkOpST0h8RHgKUTtcjFw
SV22Dt8PLTZP2lDYffnWlwV/2pfR7ZuUQ/YlLZ4tbgsFpYxk83eA9L8yXwVfahWMqeaWB/8xcBmS
7SjlouWV++O5z3U/FOEYj4IWr7OlGYFoesFtJ5KuSHOaCpDPrJDBOA5jc0c5cLkvatBIWFlX/Tvv
+FjqjBVSLv0gw+SMf+E9AtfFW6pfr0e5uW6sgl+WMsJsDZXzDEdnpkDx58W9Mbxo3XfRMJnkyjNE
72S5XUCIJOYqmYAUALGawlUMAv1QASf4HO3ki2zZOtd3sPzoEP0/AwDGMs/aGeyGW3Sq+LjETHpt
zF6O5nsHVt+HtHhoKBom1OB9UoNeqkf4EH/Fi5/+G9RNyBP6SlTb/Zbnwel+pm6vN9g8XV3m3jpT
u8nBwWuTu5vVPJbj8cEKkn/gkNmDHAX9RwjInqZPVXFmfit2fo9KzedDR+gPlt8/c6DMFKcbv1RD
yv5QqJCSNQs9QiWpdJ4Xrd0o8FFf8d6NZVhN46D5LXuuw8On7qGmjOzOIorPbLczCGT21fKDvIiV
3eYXEj1AL/muSzgMYMlkpFVmoEz+VgPkFtFaNyJoVKEts6/sSuDpVKAo3TLHw46w09NuVkiJZpQ+
mvcLVmdekjlWflprBKZKtkX0/KnggTB+yyshMOX4tk1Q5u/WOtNzI0SDzZRu3b/F3lKxOXvuqvNq
gY8dwLrqeNmCqg0u2cg/kvxL1jJl3NIU2qKwEvh0tfs0AQGfDcBbQCqNE2uwQ3ncOI/ZOO4uD9P4
jf9glmOiPzkVSAmqZXSgjeeycAym/vSXMAUunn/aLrbAQRjW4sZO+iKmeyITM7ybG9l/LeR2xWdi
n+7eDmey0V+mPJFupUnfqaSqbXwTZsosFmpDwmvPUz47tUKFjy231Ch/ZCKGxSpYleOKpQKVUGGN
lHREEsamWQuOyOnAru1Ggolak5dJn8TtCxbm4Wii0p2HQgfpd6LW4daYybzkM/8xn8YfoAxqmtVB
JQzrWgpdFL9tw1P4zdDulG+s6JrGehluK6qwnspdHzaLj7W83m0wEGXvcWYOjrLaiQsXepbEoekN
xpzGSlzgVy7XR+YQwUse6NAitTiqWT+H3ylu1cL0hy7HDJz1QVbBJOvwCcrltjJo6lfotYjAItol
XCPvoSk6LsvFK6fEYlCpSejthoVAJUk7Wrh2AQK/IV3KE6Z3SfGX3yedfAlizu4K4vEPgSoyrbdr
VnaIuKxRF9m3hlP094PQgxjljiW75obBBLQ5fHtSfncqlUF3JV9BNnuoxZpln3WcWfpxrZpw1oh5
G/Xnx9I2y5GQmCD99yaucAhY5e0XKqdaLqsCIdiRxc3qSw5nuJP5PMH744DrhX62CRiyvyqbW9JY
+tqj1hAj7nMpmwACHa3ZdEPha1UMf6wLy/0Q+qfoPg5LktBG7t891d6Bn13hsHOrqmgiTFHO7cu0
X/dQMt0T2FwQVQyKLU48bc1/lf5hE5OUH4gxWTwF8uk2dHpZLCwBV94z+D0eCOmqYL1pWhsR0+jD
AZVRSoZlHftjTcdzWQ5auy/areJSBrE5eWY8nR/jOR1m9uO2SuUmmy8op5YnVLqnLamlKw9trbaA
JbR+gM0LfUma18eMPjz/nQjFmLTsWQCCC+uoCIlFn9Dvu7M4Am9Yk469v/fnO0US9hmw1HSA7HxK
ClcpUh1N/HB8GnDYVkQUhNo4TH5xTQPw5LlEEUOS2JBfl1sdvF8bCmABFcI7cyY3rc4INkZ1ZkIG
991CTLy/48NrIJSDY8UZAYbwKyj5kv6N0P92VQqfgMSf7dRwDOgxYVIH5bblPeD0aZVXV8UkIT3I
YeTmn93GLTZPxnmQ+9Zk3hWOI2XhrLkmdU8JWxmHfu44jIjEVDNhuBThVP1njgBHrm76y1EmzQUc
uZ3D8/n4+A1OJHarN28gGFKfOJCkhSHpWhSCHYfsbqcOFLMVX7XQxhFxsXDWHGtNqGilWI3mcTZM
7FvdMy0MW1fD1EfUshEn2YhWeevU+VW7eoY6h87t44h+Sonad2eHWCd6bCjp5NjrvZW6SOdbzIq4
IgUxJSKH81u+dXBBHwyKQcnStW8PoTdD6JgPSxeHZYWZ1bW3vEBUCsgLxB5NFw4q/7PTn8t6hY+5
UznKbwOJQ4rEtk0Yr7AhHScntBrVIbDajXoGvwCy3+9sB+R1snxZey18+8jZqWC1ZTdfUWBu5Nip
+du0CajkyqPGEuk4V3BHC13F0SvMt/6IBnLWSizoRz6ajV23L8zRvy8pqVjYqZalhpdrrIH/v/zB
l5eMX4R9JcLbKVazFKr+7TwXVlbnG+0L+wRi1GbYLLkH49MSjVBV++JJXpUczHlBZ7SFUYYDe5XP
+tPM5HXVzZEB32C1YscOmV5pbxFRbC9yO6Zz8A3E9C2+OAR/oI8YnIJQf2SJeFOBZ40PaLWc7aX3
flg5GB2Y4ugsqB0YEvKTTJ97ZejfNgXfFz48qWtR5qOaMJ/RUkAUg8NOQXy6X+DAdOof4SikgI1A
06kGdGZFjmFfr+xd+7JIvJkORPKcCSDAQMEq4nvLvtOGpvQEHmRSk+394i1h8mUTi5rmH22Wlw2p
IcgcWHQVh40u5fks8GJOlWa90v0obygh7wvslu1wQZelbexuDkqo992jQ/6fQjg/FAvP265IVAGX
DRPRQs9c52kGJXs+C0/aj82ZF57vXCL+r7xLPg26CFaeWUHBWygyNvdVWciHVhh7xj1MVVw1Mx+4
XVukYinNNAqpDyMEzycwTgX5ir0PuetWATlrJMinXbsacs9DnF+La9qfuCXf5V/0BsTLQp4awsO4
qRDMV3Ow+V2v9ShjVk+JGlJ+6Mk7IdBwkIC6mkfFF2BKE+VTufYtiQP6eIm0iqVYEgouJPCJ3VYX
zJE09VNSTVdSPZXa7FqrrfbwZgo2hP+DBOdl48XRdrf3uoq8dG7Fkl7hE9F5uduuWE36X6OzLQaG
b3ZfaHrk5b+gpJ/E5wrvtiSBQE/U/27hddUSKCFinXht89FkNepes3G9iok92S/+7bUBAq1OgOK0
irejsmzkNjBWtUZS7sigkZBTueIimCe1b84K+F30nMX5WjVzbyihw2LKYxZzAI8ko9WhQEs3gBuk
CoQ0Oj0kfB33pfJ1xiw3KBHZT/WOyuzsvBbG2Gcliupu9umyJtmSejKzVvQYEFdUEtKRSWU0WK9e
1c9kHW+xtFbF9qBYcidDtCnvWJtyCZpq/hb4n752bEXOuJGDFJEgDkx0YtJaTIjE0HPjxHuayoiy
PweKFPDix9IK5jAamQDiK6CgHCRmPem0+Jef86lX9gfC9rw6bsue9x6ByVgyBhd1ypzQkg+hpF1K
yv/z8GIHsqL5dRXGuDXyv0xBoUnuOH6lscaDuxKfoBVCC075hqdTlbvmQFaLFGI9D5RFv3xOGQ1w
J+IFSKcEYHXuMFY1SAzqIVzBZvPrL30BkjqzYgCOI1EliPJIGynffVvOBzxvQgjdudQbM/RpgQOS
u4zheMcQLDdWTW+kTWy4jkhHbjEwU3q0DLiK7ZltKfpCgUldasTp58mmBUD1PCBY5NnNRSa7hcPY
oQmJNQraub48naKFBCD2wgfv9Fw2yOFhR9+mTo2zkQFpnWGJ7a4EfV/ew4yYdiNeEbAjLmhLneWm
NDlL9p1W74CbhJozhK0vsOVF4dClYMK0PRJQuq3rXRkutnsKSthompW45e2m4M3D8cpqCYBGoNmX
vhPw78GBgSeknDB/8L00qqFvS6BR+yv+fpH6xDRiU20b46BdVPGPC85q02pKvdJxH2pHURiK1cA5
tUFpaWnYpeQ7WZFmaU5/DDQaT2TkpF3QOQ7cqqWte9WC1EyqnxdwchTI3f2Ht+uYcXHktHD0lrOX
9ICousIiD1xxYQYZWNUdAkBdz6l7wPZUtargVT2hp9wzstz/69aSnuHjdyvTaKNDcjCn1DGXpGes
AJIfxD1KD9MPWb5lpLeZnOCGDrLAqoR4Htd49vbNrpFlzbOdiDHdyMuSHvhUGueLm8qmG9Vy1/QV
/EeXBqELB+C32EQ5WPU/uzE4+XS1/JBQ/QCaMOhAmVWQ0+eNsDtqdvGnb252yfAChphu/tdm7m0N
udI2ddAQrfe1THQECjKnx6VC2WP7pXA3CcnUu6HZIHPvTqnMVNZkPjFgv2/OWIuxwHrHZTaAkY1o
g1wqbdvzIq0YxeNkH4brWjk7RguwWvV3eOZaqcXfKUmY2NMNYdyzOjA+TFsHEj+sfj98a6N51gnu
9fe271FXZWIMipStFOm7ESfzbFvr0n28Ca0MvI1XhAcwTJ2AjN7Z7+EQE5GPp3g/uX+sg5mkNSAk
/597wdVs+HYhWgQ86RbZvdVi3z42qi5CDGALA0UgEkR69mgaR049D8wOADDgJd0fYyMD4WUG4zMR
18jug2O1rl/A+uU3MWLfDWgubocdn723+KjZA/nSgw/Px9UFJ2Ii3+RKu4ZOweUdUV+VMzKKn9Bo
9/avhwVNPQzXYRpupumn0aAmCC/eWQEMiecxGTjJkriZJvqQiGuaqEvkG2j5UAzSJW3+WnFfUNYm
/BtrjtRy+WUIbUF7e8YjClxMKFJbhvqB3OKPLwf3vl/n/kc94DVihbq9M21+nECaiiEQCFwQsVMh
ZEq6y2DwuFUyVcMV/7lBTa3P5sGyXUZuR9jhQ36Sp/Gy7JZoCW4ZHsX/HcK5YLkeGN4qFAyDnqVT
cKYQPoHd2Ru4xnxWo3/xHN9sGxu4lBtFM4Pkb4rjjXLcHjHzbKLA0ZRT/FHdnLXxA90NVMj2xgM6
VwaLph7QgXXAJP6ro85c9nTUvd4fjWaFfQDVU8TFhI8YyOjSWnzUy2Hefy+yep4rO8wMK4P36paN
vtOXpWpAMz8tkn96sY2wikPTZGlrBcApAcQ5VbzrCe6wCtl17v0H65qno8Pj6hKVfO3pBLyzEoiP
/uJylOz6sLicAPyOgq9nC+5tB4vJISBqiEKaQgCTWWG2S6fxr5bh6r8zwaYe1BlWuMIRUNhe6Nxb
yrVf6rQ6XwXUn3Wa6SdtMfv9oSgboKd1bYSMaeni9ilvCKvRcxDO8130Kkm3NW+9DLA6b5Kre56I
Hwl0Hdo/lbgwrLnd2+iaLCamfT94TjsBLn6k3fEvUbwkcohp731ArI70s/P57MezfAZVi6nWxD4g
MiJnyhxMsXd03EUrj9HfvF0NKTlThwXu7/A6oeTrPZtmhvnMpwcgWK3zPrvkBqVIapCalduphi/L
Fnd9M1jc9ZhbLNDluXH2ksqhUkTJcHcMj71cUCevdFJ/6ytpiYS0Ujavmqyco5E4fMCqUeLh/RAX
RHOK1Bp+40CraQ7adSx6/R2YZH3KavtAHTuFOHSaBIDhWA74XrBYyiM5Xrisjtk+3+TBVHjOxF/l
8fjFO6K7TZeS5gUbZmhFBuV0VJdtfgZOG0CUsKxdzVrqh8b6ODzsGVjLXUnGrwUr2roBRG38vlEC
5nRu4lZXi+24BmCgGeNJwYGqOR/oBmkBX1WRO4Ezf1FGKm5XPzEQWrjhKuTYxdJjMPXtl/ulU+Hi
vavCySkO+NQiX0LrkgnGgE4VNQ9To9Mow8WKbiLKAPv8KakrY5DGBPiW3F+9gD08E3ZceIhuAwd3
Uv+Mk/DtizG2h+ec6ZZLppl8aSbnb8o+KtueR7O1/J5NKXXLichvH3kDcN1RAcJKpNjrYbqJ8XuM
FGawV7d2DdYGM6zi4nnU3D0v6eX3q4OfP8od0fo0HtHNabpWSOOF4o5CH539y2wYV5rz86AJn9DD
9l/AmMzTK30WFuBCzfJxH35GUts1NRZ3YIBBqx8PWIom9dZKxS7IXaArb5f5N1rXP2xcxMs/YCr3
srh1bGqXmsx1lMdUyvpK6kvtghvx6TkXh2dLrw/NWuyhIXjJFmJsDNEu5ImLFvVWVsdG0iC1k5Ru
Y+1Ps5Q7vmSg3iPspqP+bZf00B/kydtbsWBNpZ5I2jArjop8VYQouuSap0SSoUYLJmZRkEgM4oW6
+FLKb6WRbt/WIswCTxmI8CcqJBufitqUGXdSXnanL8NTK56bAnxQOUeSFCvk6iTFeM0c39Prpf6f
0RyqT/ccDSBV6PY7i0r9AJQgBjpvoP4ORxanCfHsb8IlnbKPXPoL9jXl24IJRGkPEPDmZggHOSgQ
zE3AajranhxX1swGRHfzsqK10Gc1KXiHj0a0GHR3CletPKvmsyVy32ZwyH8G3Yv4J4BMcq+3WQfq
pipeoAfnYA+pHfkNW8p5SKMqscdx42MtWTsyZFjStwqb34LbLgzBDTNy0kUSh5RFeg9LV3jvTiGu
cPPb6/KLh3HLOhyD+cUWesfvtv0CdVWLXd373KAHYKO75YMpFO83SWSX94TbyX7YYRVLWc/s/edm
m9fYnQBxt47ms7w4eA4nnQ4+5rvcQRi4sAyB8EPBBhvhQIGgZILlzU65coyuv8litidHr8NBlEw6
rkSOIKfOyWKdveU6iEnXTaNSRbxuzYzXXMFjbz93qGNgAXDSYSDpHIXGi9BmyxsGFhcSqVKWbDZz
KNbWK1Ec2de7CEKkW7+aJQXtxLg/Hi0jmUHdS+INg2/SpzUXdh4w2R/3i7l8K0OJ67LCbVooeSoI
Ajdm5BmG4GGAi6TgY8Bn5f+AxXxTRf4LbwjtTvpzhzfem6lIef8SmvphJ5sOUz2JRfC75slLVBjh
PVAu0B2AGiXt3jGu/9biSOiR0SVRa4CMgDBC8rNY4HJ97yzAcxDerekDXxs/Vn3ru2vpgtvUmSEn
/8T6LPDX2CUF2LT9mc2jgOALB1iJFllDCFBykSitF1SRkAV/VKRh7Hmij67pv5bICKKoR4+6xUnR
jt8RIed1IRzPg+XIQZf6Q2dFHY/LusB4jXf1U9jSbWxGKnIIlkN7qGkisAEOTOOcJonQ2yXd7bSE
w0EiSP93jw3+/zCMXXItMAyOcKDuCQ7cR8Rh7q7kCGD0sn8hLqKfvnngaEvQnOSS1xcbz9xQdXnX
Jfl1mI37USMwd6ocIhzQ6EfLMPKrlR2/Qith53jczUK+LPhg4GLy9aCtRdMboN9XMajzzhshFZyb
5jt/DO8svTcOelNkEbb9Qc7VM0SrspCU71qhrSGH0Pf4M9Rc14QAi+Que+QlUgBTkY4LqOzLEwYC
l3kAOCUHJHWvgLF1UvMM4N1CE6Zz4aTzFpf68CMDffExPSvTSP5bq0wG4ymybwj9zunsnFmoYTz5
j/WNh3x2Ez/IflB3WaVOzOn9FusxFqEBA0EtNNrxysp9Srw6rsSfCkcxbpdMmUD21ShNMHNIYfmT
VudtlwQ2+pyyMoiW1+nL0KM7rVuYABLKZOO9RWpiEtoZjn7m9btq1OAo+JbNogbsOtWXFmyRKbtS
KJ+SZCRfekMbhe//K72m1KFLPItXezwcZaJWPkhdr1e7fPAH9k81xhM05RDkAxKTXYzVY5/MGirh
+VuQGanEByhOiBR626cK3vws0VeksGPKt6OlO+5WySgBq7xHKvsjSQSs/797WeZnij1U1aezLndL
cJrLV7Uyx/xLh9dgAgso90EBCVVmPiXt+9AFdUcvYxFgH8q9Z7i+Ipj7tYX7FHmM7eCKmWOK+9fJ
icS/6dyrTgNn+2ih3TEPbJQWZC5X9aSYS32NU3AobXnUc1ltHk5X3y+zrX4Q3GgcajUQsIhaUuoX
l5+X5eoETJtF07ua54nBNlhSrLDOF4h4UMPe4amI9S2NtyCqcU1RDyBgRBNuYsEAK8Jn/nokvWzb
/KKI3Hmh/JDn0hS7n8O4Gorzv5khfAQq8E85aMkWn3SLEAVjwjjskCRKJnzlTK29a2hFI3SerLk+
thT85P+0VRAC/ykNFaEE24MRo/LQ/B7e2sX98DnWcwOIXIcvZtobNHznYfSD0/+XGhEEaKKSvzel
crTcn3ZL1nKxJh/8FtjRs7hmiOn0/0Y1jN9sWWbsAxUGKQfSBbKHA98kJdhr8a2fyYjSR8CKa4V3
BqMbV7hxc53wdUzO7wqwktDBvPic4uerBdn9lqqiCmLgg03KadYmcCws8emQlYD1axOEIF+uqcmO
h9nrPh7zJSk9HEzHCsFKlENG6Ymz5JxdUBn5DzxHHzlFIskn3v29Kh0h/KE6R5V4YjaAeIVKDXiw
m7U+scT8DNotL7AjjVKx5OpZDYJCtoJkBk+MSWxBayBkMAARcLXDYTsjUkYQmPQuahJRgCyEHeed
lw+dbc/2lr2wfQANPKSXBM0qB9myX8SLSNWs1Q0jayB5OK91oT1jq4EtoFzKoJIA8+l0FuCfmgrZ
v0NislG7T+O4FP+9I+f5gLZC+VAurbq+o1S5qDsQw3vU+m0dxSvTBW6NwSMAV4XhD6nVWf1amEfT
QgDDJZMRUsvqVjJqRTGBycATkzvIwe041Z2torqhS/wYvNqWX8z0BRXl9FeCVMK2IwdneQgqGjK4
Nrz8yN6Gw+H9ORK78P9KY+OIx9LN6jHl1BoSHeE5lJDp5qPPOg6XWgJgMSF1ZWFutdV/clROonSP
yMgCeXc7e6sh2hvqEAF3m8ornSJnjJ1h9Z83ak487OI9eDLL5pojSuT/qnK5darPJAkfiVkA/qu6
mKG0T98hjpkOmV0s88oHB6v0GC4cp4lNd8cFNPYaOXdTYaryaqma3hYOZLdL7MlAdc/h4cf4j5et
S1n1/aTJRb/p4HogbBC0jPEM93gKuoF73COlkf/z4bz55FHntY+UCoMBD+Oes6a4HHAI2IuijiF9
lRW+Zhv1SAeA1XKe6EnEOrAXxcyymNzm0MVqNKPhbdXq07zqq9/UgO7a8Hag/UW5eOjzgCl5NMO8
RjqTLnrBAEv659H+XwYT5Pq2KzOYu83NAPt8qZgEI41X2ZhavMbwzTyjBwhdRQYLvIGQYjZnL/Md
sRgT0k/sjmU1cqWtNvRu3+zNsAiRVXBpbkhAyYK0pgfIU1ppsmtiiADYfF/JhBJ6e9MF5wNXeUVd
CYKAB2yDxUNHAkTJgNiaWk0i3OHFabzFb9poWEevRGkrY+4XmBBPftxwYytX4OeOKgIi5aSoysTI
hbizdowjaFXFBTCL1zpiw24nZDBEbb9r/m3899cwLCCvhKSzKpXiZvXCdmADtbPtfFJPa+yyAcRr
huYcyTQpINXROuna2JrQ0fmtQCf5hopVn+U+yA9Vv32Lhpb1FOsdNNoAzrKiWGXIeumQwYAWh/pX
0bnP4aBuSUNHc+c8rqfnuhdCKOd0Apx2Wk9Ox0wSweshKd553lUdgzDMat1X5zEgHqkoW5wkghud
1u1VDHte6DYq6a0SV8PrvDJXkGnF0LJi7A24FQgj7e1F8lwo1aCmrOY6uVJH/79bSGNCmxmBrCSr
W0asrw6wjbtDR2KCqlAQlv3v+Hql4j63L2vQ3VCZ/xDBuB459caRX2z/7KobJ9ZGj0dF8l0kBnNl
GlGcGzGmDG6DvG63TMEkqS+m7RBQkdLQnQwFmuexUp6+sW3Ci0W9W8r8yRPgI184UQsRFJc3sn4N
lkJAna6rxNG+6VfQ3FLfGnaqT2hIl85TG6ehLwpOPGji7A+YMVf9+sa7O7KXLOGz+hqrbRsFpoVg
T/Pm++i++BQvB6woyuJi/OXlOdjREBfV3mzx1pII6QX4lh0wRTANWZ6g9Tlr9vYEvSIERzTYdnrC
Pb2imaPRyFc8mMEjabhfQ3zI4/NZGeYQbB5qM4piXabKOa5kEaLc4t08MKCojxoOD/cjmY5LExVM
cGqXiVJNinxTNiVpG+2aQ2ZZT2jxdl/xFpwgD8YPZnv3CXBmIAsYxUXRIqfJedCHQNU2VUkXwZrg
8uI3CxP24OIjmUa2YA6HNrkCAWT9GZBQ660e7JZMt0AtfXYXY/9gvjXF4ZsJNrTF8nPuCWeqGTQB
X3kan4pdD4KAr9uD9mkX52sqrMSusPIsAgfxQr2oR39I3JZ0IeygQ78ijagQrBw2r/9fmpKa9Jao
vwtnTnJkms4reYRdS7pjzxldjyb6Cpk+RUE7+7Gfl7vRHCkJYDlSNUN3Ns1c3JuPinrANOBAh6iU
CVVXK+aFKPnvrI4AfaLDXOIBxdXPg5ZrSMeDfR89QqeAK2JhSPJ0o3cLKtpEnnk2uaDUwebAhujA
BWmFVS8B0eUyQRoBH9C5yUW15LLKPPHWJaqQBAuFzYS01656MGZaTIz/OemidAxg5yV1JWYAoJKV
wab0SxGMh7DV8AAXBD3TKOp8zyxHJaTE55ENp2EuzTOGuGfhfOb5FDgxasFNiy4VdK/FiWqQ82P4
lsrNca7AYzFBIM7RzERQPkiq1XnJYINQ6AsO2O0KICk4hhzP6NUnsv9iiE21ZvzR/wZX0aX8bLAm
9loLU4ztIRsD7TBHMJ5aYaXYhYHOYVd+SCz7uLrd4YiO6tE9O2nGIAkMMN1253ELmQLdFZJR0j4g
q3JIO8nCMoknFsa+2735rRaXe/vpwOYwlFA3wpzwGZqRG3j3sFgraaNxeTyFWzOdSMAhTaBJ1yuC
GYU5bnOuHhJxp4E6JV7wQ/ebdqULqAP80JWuBqs2EpP+t/QvdDO3rSpJgC10em555NOi1JV3yFkM
z2lqDMf3NHPtvrARr21wgoNzCMYQfRmdH7u9jjGVCPF14vABlL7CazthZbXDVIhi7vBeAtzd4+cB
VrfhrGPxcIOUxTWxlDkyM76cc8I3HL2QIKthqqwD3958eDaDDOqpRZBlj09fhzG743qVmkXql465
5z3wWzkrxg7n1dsn0y3dpUaVXqIzvVskc8oCcwEdgWpHHF9vs8SUs3Qe16z01Y400bQBagtYWjeC
tnjgpUgl4a5ol5krQ1gokoDU+bF6wpP0HJW2V4LBt5d7NrxHpKIG7VrlYYmlQHXFjq1hP+AgRxVf
AByqBeM/JSs7QOziQYj9Db/OBgT58Vg4orINCSSNc4qH9d+p6dyjusph/OwdG8o/69zaAEhD2kNM
cLrw1EYO/wFTtn9gdxTbx+yDsKEFiPUlb5u3WuwHAuxjylD+v2565/avZRyqNqGlFhp9BDuYfvyo
JEtOXLB+yu3Jxzy0LAXwEv7BRuD3DjGynnIJ1vV24mX0HOZ8/vI0ImUMO/Kv693ALSzOa+t8PAtb
faJJrl2uknp/tFKOk3uoy6FwoXnPRyVjvQNwdlTf+n6bekWKIRdZ9lA2LqUxEkRfi9VU/V+qOPgw
gOkzE/NvwiuAI2q4mp1Vk0kY+iiVz/6c08vsXoTJmsZXhy2Wi0qDTAT2oDtNwgr5hAB787/zv3+1
tsGGoAp2Oq83R26QgiAKTTm1gCwqjL8TEBBrJT1ZRM0aaS7gZWiWdSedLtu1ESfcj65jnNZnezUj
d+PpS7e0X0iOBVE38LgrZRwqapJ0VRlXwaIiOeLF6gVAy5JpQg0R+EP2dnMa1rV5G82DKdvA/Omk
TGLIYUYvUChGfwew7z/gc7KKyj37J6xZYNpKiHTU44PTn6kYbsRd9egFxFholZdmwjl1ZyzvUKko
lxKbGzLLTwNo2pVfORQs69qbhw0B36LTrHVjoUGrU4M3Mo2bimYp6lCt10E5aq76WwbdPhAFRjbS
TfpEpwR12SHmYIOC9L+AtgTi/HQjxXoCwt6QN0DFiDBqB45FL5SkTUWFYqpE6LBJEXNUXA4N+hSv
fPgUDDuVrcA82BGnil3E7TDZ9gg6qG0ZLmUUiAg5dkgRRHfjV/6vi05SFXYT+HDSCEscSR2uq6wT
IMuennCE+jrCIB/Yzipb+m/xqOW3PQ62OT53XyO+ToyyirqlvbW8zZ1fl3bASN+wHPR54S51Pbws
E1oWJpH0qY9fnwkwkk1+dNanCucnYU6cxYeFPlyFvQZHMUfRNDkv0flmMeTujUxBFJ0ffhAaZQoW
ZlrxBPnZm73jz6xM4WoZlS+uex3kjIRJA/QY7UgWVPOsMPAma34QIkg7FwEu7cCT0YXZxzx5TIpq
sDMdTj6oFIb32E/IEt0QSCNfWGKBaJKDHGjjLmux1deZfPZQVVaTK04QtnpFaHDOPLR6WOY0Llsv
xknTDmGXyFCo9SPNSO/W+/ioyayFVM2Il4KnFg337aAfyWLvtNy+QsrJ+KtEkATlPoqThHfoBdva
hjwkw9G2AbfWdMugzgE49E1QnqOeWPxt7gB5NwSOmwQzQ251QJv2N3ORTpkzV60z0LTZD3u84XEt
byDhjY6fcz6Dzzm7B5NcDAO2SAMnV/Z9H2hIFMo4PW29BBCQY/9rNNvD6HnfItNDOcyfKe9mK+Jg
dqmB+Iy2ZbjzMy9MRuKr1ZG92sZyq4xpK/nRUlOOrop//yiscrwfvC4cC+vsABf99WsltmOuxFmB
WCf9R96fgkpT9uruI4LDrxvZ81QNSTK6rH5ltVcOXTi0drLcKFnlqSpUDxcLSHKlGwbZIZKjn1BI
E46WGSNoMqMYYcwxLRoM77UzlhQzlfrjYfZho0oEwEItqvYj89Oas/32yVjSazckkICGMwSDNF+k
4GgJ+mzZwHhnTrJPb7xWlibTJp5Fg216JLw/MgnHu/oRcy63TxP4gEXtA/orBcIJqwiIcUmVDmSU
6v9CW7vILb7tp11j2Q71NzKNo2hjIEAXboFR61Q4BEBZYNKt/8bNVKwm6i77J1zgXei8j7+7Q2TX
sWan2u3mQ4xqwrAifrVA1SH8gfbJuxjYvUrq1lOyYxr8HNP8O6mMhz9AfbYtDPILIjKFpGWP80D4
acxiXfTMbuc86lDi4Q0Zw+hC/HOkAV477SoiE965f/qmv5DZFggTMS0C3943zqPkpHBaJSS8e9px
Hc5JdsL49KfNl0LhNWlfFBWR/K/W+XnFOzxCrgioLIwry4g6xXdGei0HjuM8iL/ETafk7jsttTbM
1HFGh93Zmorgr/utwoN5bSOo9ZtrjkBBSdq3Z+zBxRe5wqLbkl8eQenD34i9L0mT9+NVqXuCECXX
jsY6aivvxPbZWqNJzbs7MWWS8mi1Rkxiu7ayLfP4bxXk+nGlBImaMxKAgNiTCNglsGlnWjKltbR2
x+AVxaj8NPaMKNKpSY7LXIVPvDaNmUTPNf9LX0DVkYz2/X4xdD9cm7KaH4fNxGmpxmnZNCC37yAB
sgmpRygaGUTSPp+LCx0/iX6cYLmytVBO+1+6TBLJ/Lyv9xo8Nd9Brl5XrR4Mh/gChHv8s4cxFRcj
DbhqPcI+BYMtt8NY3c+wXJFlfcEZ99WMCZfO9GQ/OLbrQr0pR5whoBaZE590NtSZwwK3yr2ZGBfk
tcdB0eG9VU4oXGSHdJMCKGS67J+LzeAbm7HYzsZ5L5593/IaTQze824GOAnlicLP+Xm5hFX0+/f2
j0MBmJL+nz3NboXxTVTS+NmbqTW8Vy9HXrgKCaeVQQJU/7FDtOvzYPB67k7l1ZEcB/nVbpTSljTJ
CIdQAL9V4Pr1ogH59O8aTlGVctrS4kbXfkXlrvRiHT2FLsIeweAIgjN+z6JiF4Gr0fW7KZITnkyx
sDZiKzYbVE7ynEkqX3TRssegNwzU7c/lpDP2+v4kpjFIUbyyEOwICYB9mJDLzWodstwWwWjILQat
0dY1lw+6pfy22jTDO10O/2QR3KH1infXnvJ0B3DbbU/seyAgPrRtTPSKTs7a+Fwknbm4VhF6hFCC
mqz0A0UG31Nh6++O2VIJIumv2wAv4lvR1T3MEQUZv1tLtpuJTgzQI7RTWbjelOuBmCDWEyizBFUQ
RvMRptQ6TEHC8Z7B2HZ9UIgvsdHOEmtxwLa+cIZH9J5W4uy8/yztYX074VNwxwYNwry3CeYJvAiF
gqy08YeaRGr2MvOqiSb2upEvrW+b16r+fK7tAOW+1o/botrBTx93/Pg/D+6CZq/w3P1sbBbOEMuR
ThgID+c/nTgbJYfM4Gc1PD6lwT4y1zZA1HfMpZ5l5FWF1uYURR9hLWvPkxPk0X1cQnqPxV7GLRl3
zK+ZOTzo2R56QpC3/IkoeLD0B6nffxxLISl6g5R9PqIaAjXMcyUAXjrQEJazDm2KPfqgh9GULCHd
lRGt/skcfTnaT7BVZKbhKZHwIueFhlCrKPbAeq+ZouTZMBEH7Owv1L4vnk0fgstKL2k3bKHbxMtP
OLexciTCPsv5KrGwEN1607bVghQKF31IHfX/NYY553mO/TsTJnkIPMAGCXPyAWsi57n8q8I9X2dA
L/GUkpi58y+dDeW8dntPuFNuK4lVGbUCWiGMOS8Q3sRBYi0Jrds+u0QEzAulDTQshe/gZYovhuZ1
VncWD1qb0NjQopf+6i92hjo8TEyGIhrodisg33fkhiY8b7JqIjKbzaoAWHKEt6aM0DIr554/QRYR
gVeCPae3ZXAP9jKqBqxvTc53GkckfUTUtFbmP2FzhqRxkqyIbUmI0nkU1yd/GGfId5J7hYuvCckw
xHB+OVeCnfxfbwfEWCwzIsMb5qLu4T8u7Kodc3V22LgwPvuyXQGmY6I1W3tT7dNGG+VoG0m1tBiK
gCL3CjWPqBX63qoO8zoSWDceWrmuKlhoB6XxPR+Yo+GIsJWTLOx9LQhNfDS3HWYKM7ICoy3QwrNW
0zxCaVLDJNy/5K42+iTRK3/394m2znzom2DuW7hKpz4EIxGFGlpV4IID4S/73MmMqQ5y2WmesFKU
VcFanWs8ZjPcs/qDAggt/Csxraq7X+bNj2GtMXFSb8+PZraAh49wFx7xl6h91AYT2JVA5BuQsR/Z
ccJpaJ3RwZ7U7wxmKGrzOFqaYr8IbVd9EhIh+Watyk1ZOm9FY+3dBlG8MvBS73aGvrDy0JiOdzhq
YWstL7toak+QBNkYrvm0IwjOGjq/WCcC7lshE4kqtHrLe9Vz0moOYeoJoCa2DYHzOrkphrY6CO4l
g3ThOpYrSznvpIGqwvRn3v7flrta7JwuosjuMEIeJwdRKwazznMH/8i3j3nMDANZH6PZTZGzEDBg
wHTSLifOsgp1DQoGrJ8u0EzgAD6rRx9RzEvzY7PAvbE3nb/gKuuq54o+Mz5+RtTVy1PY9xc5+yVP
9x0byF1YJqwl5o0ZZo8zGFaiYWXZqdlwB4IMHXKwmGFO07PNc9Ipfk0aJcPmsppKt1nKOP5A24Z6
EyAuJx3DCnvfukr+95iEP2QQHsCJNmjUzdxqdMHoUEZjaeM+I9KuR+gI1rXid8PI1gS6Oi2svykU
b74G5Gq4mHqS3vORamS5KkAzZBU6YFXEtSOTb+NSLF3nYdLSN+waIwW4fuK5PVPm5Rz/NFFB2l3H
rNFV3xP6f/9RI3/+LvcDRyxKZhH9wMkIBtn51N1R6XWMU+i4Szkac8kgEMAWBOHVyKkfbg+Xl0e9
ZI77N250qO+4UDKTzD7dIGOkK/tSfTiV4mGT4lFtc/GxW61iKkuoqvU19Eqe0eOIPqjg7QzSIUo+
u4bL4NXTmeJIidaLH0Q6hlldjbx24SRrDu78+4tEAAGfywEbQ8ZxUOyvwSaNEEQkFb5PwIPfrU3E
076qlVE5fgMU4Vm55eavevMauaogT75qo5mLfyB0B6nALmg+3RZfODjP4y9EQ8Rl3MgVvCsO7ndA
pgLEWzK3MkZx/kxDKqCGoEnBmTDhaGMcoIv1YoyLu6h3Ia6pHQjAvCYoaMBB6bQV6nOJCnh6WlQv
3Nsk7Vmn6f4HhHvWXblbX/DCZXZgvDaHrdmMFoWtNjiNAsfGz1zIMr+Kwsz2f4DJiz7d7lYZ0tLE
CzBUlPUT/KZPvRUzYITNJZjWQHg2QqO2HZX2PvJQkoKyP46JATh6BRT7rcymkz5x4tASjxgEIY6B
1zngf4u/jeuC8EGUu7NdPVHFPXqQNGcJFkYwt8CaBSyzZQzM2/YO6Oxq3awCJeXAzPYH3iJBlbtJ
+2czPWy/8y3gJa9KWxNRSafyh577ojcijvXnt5xSaGRpQhv4sarIZ8X+XQ1mNT3z9mMMDxM6DD27
D/oXJu/s40cwyFPBffJWFeF9nLYjQh2L1WiTJhJHox5JZVm3nw3825nlZpLnPBlAysUybOKhM8Hu
E6F3GBl2qbMM+i/Yd0I/mRx1PydsJ521oplvynYBQ9ZfO6l0fcBcVdX46kLMMyJNOLmrGRK8S2vG
VnihSO7k1r52uZzuY2tmsdQk3AdXjS3ux2G8aRLFU92n1ym+a7cj2HtS7Oo+XngCA08oqKwwFG/6
U6apIPd1BO83pQOib0G0lY2bmjHKcEQm/MtdWoqfIheL+5OQgo1Tcw9FDn7NkjkgHr2FnXRvN5Wd
il+Gc1i5UGwA2UDlXywmBTPANymaTgvy6GTN4XxgEIOfT/FLWqsJojs7e6laJiIfkrKZg/HgRhIY
qjqyk2rkBnpjuxUWaT6yiX7V+u2D03S7LvxPfxFERXS+KEMYvBnjemQHf+2xa/GADXoe6bPo0W1b
g8PyF5+A9FoI79OK9/BkvGe6iIkisQumc/aWKsx21+ZQacrYtJM6u4fSBmwoCP13O8KRob0ssWmY
Q06zIZL8pJvGXj9rfUH/8I0IExkekhfHLiMOuzTxCCuAnS4XLzSNDSXkef0q/kQiQbakyr1S4+v+
lsjoPczJSyT4bO5PjaHxo0EPlx5GTLHftv7/LGjSnCuTud0Su8P3t+xLOeboxkwA8UbGyaKyP65u
JLLOcm2sH4Teby5qWPBkmKK3qMgoiS22FfxcPQ5WMFbxs3xENjEP4LO/8bu6XOttOMCMZkOkPBXA
1RfSg82ETUIUtlZGhAUV6PkSgXMAhGie/aoMMKOydIZXyGeXzAcn6HUsEzxoHjCckbhJooZijiHF
3WW8Xe+QWoQbqkSCP8tRjJmdA/5MNCyYpSxUdLXyF7AAqBECRQbAwGMMEFKe8ZmK7S1erROyG+nb
JNmoGMmkX4u7yYQ6/VZAXucjCVMTIVD0rCDgZ6aZCHaGT8Sy+xVLdVi7WZC8P94cvwtBAhmZkNnM
WOCQcpScpkIiA0LA2+BvdlIGPD+8g5HSqWrt4SiShjoVyJoyFdc1Vd0BVy1ws8HHJ8P6mcyg3Pye
lSHYbffjYXF7qD/K7sWs99HyHQN8CEIUxbL7o4Z6ogDLeBiXKg6AHjZFHNDX5ylUGAh2+tJiI2+X
poFDgYaAEf6q278x91DphdWdKJ7+4JKXMmP87vEu6CnjpznUSUocd4SBF32P/ph1R1SjHGKS7XYC
GpAtsIEydUnnOBliG9XgIoRH+lDYFUusoHQzRN2zml8utiMNq4CuxSD4muBLQcGKw/NpbfPHCUCl
YpGsyeYMI7mhiyLWsMjJayJApmNI2o3Hvpx1n3kJ2m11wboQAbdQqgz8TCa8DJNtXwF51H+xF7qE
1goy5ffGw3JxWsb9l8Mg7xzmRzjybOHyz+gHDLoOx6uS/cBnLXsP+veR6Hd67ntMTGMVoRQXqzFw
kzss/aItf9vwdz/U1W6IiH5ay6Iiv+4NB6p8vFCMEKJXNUqNceUfi/Hn+f7Tyv0/fLAkECSa1O9B
FUFegmIQMiaMWnq614Ok8TlFYITXgYR1HYvQex2razAvlSkJ+OxAoQ0iVOUvuuBhGjvg7HD1xHh4
TSM3aBfvNo9ZZLXgfZoaAQ6HFKq0GoztttMrGC7LttmNxjQQy51fZEwS5jX/8lFsosPcI2P7nuN0
Cq9fLP7EBt/atEkFb35dlBHAWoiNREBl8I0AOmYS91YU0ETweCkl1MgYGJyia7NK9anXJrQT4hc2
5mj8xqOvGVMVp+F0+NXSn0C2qYI0hAhCwxTRkOk4FX2kP7yJxM+S4pk/REzMouWPUfkEyD98xZj2
E0CzbXX6ZvFoO1rpFrJQf8hViRaOczIZ7Af7PloegrlDYNVk6BiGeNg08y5BgDZnuzcKmmN43whB
uge6DtYCs6UO8POv1Jy/dLU+QOdc0bArWQOfh5SQNZGsP0JPJE0KL+2e/q0azNHG51jORH2EElgl
Dr1p/AM8ls5AoovjBrA32NQqYd9TC/e7OnwZGJn1sDQIEbJbquRBtSp1zrLxERRdDoZKK0zItEl2
Q29G3z2sA8c2IioOP3YMTDuNR2iJ+wKTDesilEpPYAGQMOnjik7EhYtOlGXAFiytDonWAx8Nenez
xOkcmtcb9DKf5/jC8TKRHJAPc2Idw2m33i88s5/h3pxvAb4JF3q/Gnd2kwTGv0BgAmyrKNLx9S3Q
ioRLvnM2KER89jRTZw6xsH5H56PnLv4qGeF++lynfpqNvpe0j0auZpYBl910F3BfdCKtZBg1hIA5
n75sR4nQS671cD1E+NznNv0j1nM85wswYiiT/Ox4TCP7SmxZplC/JiE2tJJ6uuEwf/TW5VtJuy9M
3bx5YdlpJtP8n39QZzx684wOQPisVYdWHgxA5zi5RfmvU4wc1rjpvIXhAGD9uhbapZESHoLbS3/d
mJ3OJbrmUV8U/KD5R05DvpjxppXAkSJUqpEZnNF/VtEZPYFosexRcqthc/EtfEvHoooDLUs3eOM3
nzrr8dOMFtSOu8mNTnb/80q/dL+YcBiA8qWcz+K0RzPPlHdWcnoZ2nV2VDP0u+ACp9FNP15GQIjw
vLmjVBhsEDYYoNK0l9ie1WZgBD3rKLb8Cinc0o/fSU+v3vJ4h59BJS6haxF+jFlXDbsw9/42xAt1
IQ12kh3xZaKo+KPXmOhyuQqOUaaxFVsxIyLXaJULvdrsfeRWIayCrlb8Ip4sv7CWx2mZSeZW3kfB
Z5t0g0gBIACycKTBBt0IO2GFRvdnV6dkkjAYx6AivMu+451TGGXE8xm6yNYRpLLnDKjbZLxJow2I
o+TDpWoNejW3gdx5yiq3DEtNnDLMf5j6d+Dz6QWgKb9zWjeriPABTtbyRpZV7owHCthWepb055XN
r0vCnIx4KxLTdEys+2AYj+DHoR+deLde/VqvBi4uO5qDk+hbJng3aEI8+prTUrBigPZvlkKM8WG+
SlGcExaZTlZ09OKGWE0eWZNYZFlGe2lEYY6kplSwQvTPUP1YJeGAnhftJpabqNODjWuwBr3aeXQF
2tbzGazsK+qPz0ZohbQnTEVUmmi/a7uUu6sdV3Iv0ukMk7gxpHdh7my5l2XiRjCkb8ctjBxrFbkA
53GEnO5MNvMDZdedngkK/ssv2n0ekAZEaehuTO0qRMHB4iRLiqNVQj9geQ725++MdiycPTe6R2PH
cidUQhr/BjlbmStXlZCHVROgMfVDAJ+6UfC01h6cteJ6kvAKXkv6ZB5Z08COzZ4ZxY5+RXx80o1y
2SyTYILoHiT1hvd6C7G0qjjHpWfK0KI9UqnR2qc2sY96I2jiM979/t0UP5IULo/aH3Cji4k+x31I
8Q4M01GFnYSX8ShJqcfIyiENxLeDdXTw4eZc0jNOL27jrvk+dw82qzzrqilc42es9r7yBFSgJtv0
W7X3/EjIUpqI4u23yCsUDjRG9nFIwo8hF3KNnOX2Vku0e5ePe2t4f6C2dqEsGZCeCGq1MNVGTGtQ
TgpsAn7CXNx+TAJYqsQk7AD5cBdp6ZynVsQOXAUphXtqwEyUafpa7clF4lXJpiD/4KI1ssFhuthj
xPqDzlGhO3F7vIeKG0FrEI3xiJh2tYiFzc3IeU8ll6QZXGvtShIv3LlEFX+/P04JRR/9moAJol8O
zZIX4tG4equpk5WQfpfD5LDEi6FoHvo0Mg0IhN11DYJ5/EdILFFCly7KrhQfxDHH8YVNmXw8Em6M
k/0iUNHhwuVwNGcyR1MwwDxhB6PAMyx5ok7ndfSmUKPepG4Sv0cd9THb4z1g/dFSNz3EGNd8smkF
JQrstl5rlq3abwfihTitCst+DIfuNjOR0atf2FxwhdZc/YppkSXMYAOmOP4mzUn+ylCDzolA265p
aca8dW/SCbU7Xe5jAQjHyztEgHpsEci6f7K3Lll4Csc1+RqC7+7uu1eGB7WyQzsl1mMRj4nCq+wW
4160gbYCH64Z2ZsN2po3JJXektd6dpS4wAAnq6wzZ0apVWFCZFgf6NyrOqDTUk5jQ8hDaEuob7Kw
gFIbHk8nxX80KJucpbPkoFGAIvMKMuVd6zj7Bu38g/bNSyt1F1Z3tzsLu6D2NHNnVh/rzD6qdpCJ
bQYObnSCsTtKT0w0AfmCwt3JXyzUBdNIUwJiwdzq/SCb5ZAS0Ntl8vGTIAyKJcYgaU4lDAxAWxFR
9qfNBSlp/7iipGbCURdlZZRAdHHndC3OM7n6gfxFZS5teEkm02swTuhbMqjoPQenqJNbEYQ43L9/
X/m8YzxPMWVFg6rsy4LMzogePXrQ4u7G6gKoOv7LMODQPay4f3Lt3L3J0VsRNO+lysJnGl1PRXsr
537caLiVEzPkllwffOpi+MY/0VZGd2md2l6mg4bNjEhekkFku2qNUTMvTjjNEky9tCbZtNGKmH8w
ORy4Y92fjoBN/IYNp5hSWjmWFbvtscB9D4KZ9Vi/CFX2vUkQU0/f68m+CV/4L3wXg61YMjMGN9ww
lEj5JF8xyj/66t2KtA8CIWhDUnSbb/8Whw73mKOMAX/z0eFKXqhN0WHPZz/URv/laWJLeRccaWGD
MySzRkYu13P0dSMz87BtlBfkZNUnLjO0YSgukGf9fAPCcxX/H/Nil8f5PjXNR55DFozdaLwQnNxi
ZAl0XoM0CguDYHDsD4eocBP1CgTlLxE7893kdnozbn0KxWx6ldnoopMOEaUN/MeAVyKJulVVoDq7
Qj4JRfvbadatzEgzwsB+T11FV+qmNvGdcwIgDqgpp5Opic1HJQO9WKvaT1NxPprYgoD0/PO5WZhj
sWx7LeLQ5wShyUXLJJ5874JEzotdwU3GbhGMWpu4kygvVuqN3VJ2so2DmRLKJhI1Qg4GW9DveQEz
UgeLYsUHFt6w30g9McRgRNKAvFarmLrBLOGnEXfExAMhYVCMDtdO2HCROKdkIbDrXMLMDwnr/VHM
AQeqRbV0coi5Ve4E6wV0n8GLdLMyaTipRf8PWpv6Ye+M2mUDvruk8nuDmwI3LmyCU5zPCpepxLXJ
NrPRL5FueZtGWcro/nN7zOhBigS6pcSrW+d6zNGQcoIgxjNqzI1pqUGdo2pewdkVzZDuAPvz5kco
LQZHOQUmp5vmGaNTo6bcl+Pqb+DImPCUVFhEYWeqsFeoj41+iQBsly1YvVZwT60PTkCH1iuqxgQ2
R9mUwDDNjqQbUqfiNwVJYBcOgY1I88vZ2r2kUJ6eqDOPjGlSmCk1fHYnDk02lK5Y4vpc7Bg4TV5W
g4Hh7AZM41qoGNwYPLmCcNZgCuFqDnTgGW7UQqeV3nkTu46HvsaZJ8iWG8twa1N+L3pYYKtF17X7
VWLB0po/cWYuHvWObYbVjNsylnu/eJ7Jg2HsbE/OOCE8CaX3MNqPW+rdN+EaoEQNQ6TszImJFxal
p8Vwtk0raLkaoIcxaY29S8nBkpZwSgTvwVgBubrGxqlRmfp6QzypB/FfauhonUTTkPeR/fLKdVqu
+W4eWyd8rTXIqiXy6flBToMr3xw/QiM3gX4gLIbruHkEPwKz6YaQF9cpolbQYxXaeO7DnMyZKC5x
k3RDOnJ9z+zbjKjYyNmZPE6m/BXtgilLVxFgpN28Pg8TAMHat1vF++XuqR8Cgtl10IgZ0L9gqgqN
TMtRsVEY1ltzMw+U85jAmRueqnEnmGqHqxwMsXSN3Ewg7l9b1izEALWyXR5l9OlOk0yHkYEJAtuA
Roqk3UNO4qmHzOQ0VpGfY2aja2bfkznuMayrtRTt5JXZ/G7xbXlUcQveiirDakniMnMPdgUlJMP4
p7fynbpf+met0oJ1voZ8QGlCpJy1tYIlTVbxZbYNKzehTcJqUrorhUBGuH3K6U2dyg2lUxBs0MFW
bfFXyij/EzjSIXv83xOpnGVOTwqG4oe0Zv8f1dl9nqe3uYB7UcEP/+NWtQ1T6n6Qb4Oy6l2JITV9
dDCSKLRr/GNuW21GOiIOCTJx7Ppx2RI5A0DF8ulYKv/tg8oIKHTFwIFawK5/999ZQgLGDrZitkrr
/aKJuQmc5t5UIwQlH/mfL51VUa0i4HRLZfPs+ikkHVTeOI552G0rP4C8icuIo8W1IlZjHW/rW0kv
HfIe9N5YiyRQFY3JxTu6CA9giQqAEpwijbNMKT6xZIF9Tf28YaSUzq2ybhMHeOPVQQBaF188P17D
w0ZNchLtgWXujhndf01I37PHX/CXDJzhtWvJKDIAl36AeywL0Q7OMvBmpxWdnLNDu0FGj3NU23Ms
YHS1jt0PA/LFZDYuInsz9M7EnhiI6mkY9At9m0Kb+KGk4nWbSyHxHGMJrrXClNbyC6mRFChxpM4u
vktXz5alN4W+/WrUdV0JYd7lIsA1gBVJBd84EmgIlGbpqos4D0PEadlpHnI4l3Qoh5qiWokLEYyx
nHdPybIGc8eGUGsLXgJIiMKB8UKptR96GdenqKPT8WhwG+8xm4bKE53xF4YsEo1RBR9WxLJemguu
BZ889fQ/pITmiifs1u4DC80Lhe/MAbB+nW2Oq7EnnKAN9arW7z7nJzuUNb9vez47Wp4hoWTFqQm0
01GClsVVC+tWOtR9/fLXoJG5EHnal9nQeLz/n7g+U+M+UXr9hN4FtoP+4MswDlvdnvL06QbOt+hQ
GOmMfqwiGwAqrzqqDvitequVwY1S5J/ULgHx7jUKk1rTGbecQRkEIGFJjQN22v811c96B7T96IsN
ktWR+xG3RQOObt/IJW3wdFfUaOajHFloPH9F9zR/6bnELqR1Q0SxcEYhilP+bimhZA7ehDtgYJpS
bLgNX73pXUiaFvy6lR2PntFfRnamemYu2F4APL/9Ykp+G4Jzdj2HsWCldjFAN2yndDS4QFcz95kz
hx14o5mSB5h2sST1Ye1rOvPY1BtERHi8L7l6LjK6+LzD1bpjZwYS8rSg4fJ0woYDM+Iwdzd6/03H
vw2pKdTNjHZ1ERIi31cPWszZvSspN20wNmlpeMnRTpfD3elEIT0zj0trsnu6uG+8DQG3fO+P82bj
nJJfrmgkAkkeCVQzozvwx3wuUOkdIZk3Dt29jdP/Ylm0JjUu2i/gTAQwvuUSphEUX84fnNH/H2SE
/1m29BlK/WvUGrZFr9v+fbLDG0ezXkUm0qGXrJ8NMTD34yQmVcy9GOVy4PoiV8b+co98kJ7UbK+Q
Ve3gnOx1zeTUz+8lDvbwzQJlMiB2Q1HL4IedDoIGsFqDYQRuTyc6C3Ft1mC4abj3VaIfoY8FMV9N
c9aFzRAQJc358AJ79/0VCZ6wXLAzabXVB/wJPE64XAmDmWU5RNIS2jbcVKBLXi+OHI6PMX9MiwvR
M1iXp3ZKcNwITOU9Vj2bo2jR/uTl+AIIDmfGtYJdUZa3w1F+olq3PLq3NCT6mxhhbhcdA+cARgNq
vRR0ZQ15S/APdP54rM7pd0C/u2jtDun1ryDUhnWTmvcKMcjP9flzlijARXoTuLQ0JkteQoWiOB5G
8Yj8+vh6+rlLhq9o0IGYYXvBBClrXeE9mcxTu6Ej5ceV4rQF6lD5XTNYiQZNpA0uQSJN9lcBwhzy
aebGTgjgX+iS0rY0IHV6Er5zu2B5O0Tp9ppVNKl5fEkwhFpRIK2ej7ecuWzMzcO3PS/UBW02iJdl
lPS2K929ZH+N37aEXtstQTRPTIfHvlfCID03jqvwti3o4bblD0aOBX5eLVyKhg7LJ6gQ7aFR54Q1
hl65vmoWX2zA4I4hckp1RrIjWVoby2K97dfxdQlsxHIfRD+Vyt78rTiC4LzBEgPCTfadtj5iWuDt
MDShrkUGtt4pLRAEqnOcIpB2sLnz/dVkVptASb+fCrs4AcAG2DuN5YQ6ZCus3uFBXhIVRKgm0cxu
MMbRBzjL2xxChnmEkoHNfYoC0t9zyXHRKvLRO6qHsVBQIU9uaMXC7eZ7tdMBamUh0vmFShnuViY9
hz704eID9FBdXCSTUqCvFvu4ZmZCOADL3jr1kgvKRFxnRDGLddIMewHBNPNc8ww6ZpMegQhNVcNp
vskRdVjqmy3WSlN7oQVAOha7x/6J9yUbkBmPTwqrlRGKv8qJnqCsTyKicJJXklYIAhqNqajcCH92
Ez72rTFbu18idxRIpsCPzMrwq3MyuJZn4B8FG6yX7assHpyJnvggsfksc8g5HWrb3/YaGVPsHLKN
KEXzx3td8LirgE2Q4xgb+27CxNFnjT96FTc3Y7sNhRvxiBs7Uk+uQRMOoRUBRzHhdT3pug5tyEAe
xQ9sI3wYt2OdtcxkAWpu7lYydAL+QwD5EX/KmdgiKmktzHMrXBLjmctSkgIkH3fe9BaQlzvaqjbu
OFkbZZZ+IcYMVpUkkE6d3nMa86XnloJA0eOyqEp7MMufGIzLi//v5VxRdiATTzeKlc2VsqfOixlS
vXXfGXJz6z1Qc2WWrtx6aFWjGkq5bY5VrrEd+inH8939+DaHnuzqF+Mi7oGPcjYsV8aqlG6SNpMJ
wqvN0OX4LyLzOydf65HntWZRiTQpgxKBtG3O4D3keG45Ll0bkqDFB3fLxtHHWEmfCKsSXmXBymY6
MuIEa0q0MOr2szyLv4H2fVjIe9dezzih/9jz8tII1wMk9iJ+ITxpXfp/pk4RT21H48Yuct1sIDBG
fz9T5PESU+RTnT+D2wsFyroQR+YcwigxvGEq9A+UVXBIOr7Cp7RYxQ+3x9dEB/aJ9N9e4RX6tRWr
EeLyioVMFKdaudfKIPPU/5bq4M0K+byWdneAmShpOUa2HIELOL9o97xY/ukhKTpp8Vw9bX4MTkZD
BH0R0RgDQ/+XMnzReJyFgbE+UzFhUAF1TWJJtZPlLKmuzVlq5uZ7rNthIGJT1TKU+e7WOTDeaj09
9OD/KCwVCT8z5n6IiP0amH8DAWeOcytkhLFu6z2Jnn+YI2QeYqlZhg9elQnzlWGt9tdSsl2TVDSq
Ms1S4WWIa01nDvMXPm4QumXpSGxlqhyH8Xk4hNvTz70z7/kG+S0zM84SH3NM9PGeH6V2Ht03mtPO
tHfaI6/ryGxA8t1jM3Wm0oDsRrkAkKL6Zvi7TOpfFDqWR5DwrUse3IcqnCgbGx5XUs7aGlb/HBPm
RNpSnXGMny9RVRBD4GrtcIwRFxJlwbxV3lpRsaJXW4DWPh/KLJqg4X8jNIErADic85/AyEu5alL3
ZkBu3V9RGpj74Du/mYzxQ5BHbGwwdvLdtJq/aY4GI8xtNAFSmUSnOVUIuTRDIGgc1HYi/bWCZIxz
OmOQaAt5ol7dgDsmBwyrux1BK7c4W2z3J08Ui+mDKwfsky8m/Q+yLN9alssGXjg8TWXPZWmtzmJY
1sw/2zvZSkBmT7674j1DaCv9HDvtpaNdmH6fr6lMatpgJ78jklWtNQdtS4Av4frRc8LcCxVyLcX+
Hb28Ppgu3c3hxSIOiElMxBGxOjem87eFkTVbAQrcoSgwPcH8v+dt9iPjH9NnIprWLdBl7+i6kw48
OShsOijj98V5Ksymw+flz7sS850GgZN1dO+9Bqs44KcqMuOHgVPd/ZoBYdOePCat/vXKdrDP21hB
BnEjt0m+Rxly2f2X6HuRkRluvg8Df2OxUBBqqHqxI6YIgc7I+GH9yTvn/iofzfVcKIPGO83k9PUs
OnXgDVtu1btdt925k5vX9JJcmdHS1K85fXhFKQ9UMZ6FJWBGlsx4owRt2bYlxuMjIgjofQfelWxY
Lnhes1vRM1tS+RB84bL50kSA54Q32BugSZULujvQLKyuCO6NnbPdM3kKDyV96oxPeOZv6Si1hKW/
IN45d4rCZ2Ac+5lSbJ86Z+RPkZ7JMFrkE9UvYvO+ZWZ2GNAmziyuh1yK91aHmmDgtJwfI2o57KF/
KWDgk+lBKQdlFE4Vc1Z7jDjtYDF6lH3LAYpenbvrumflD1DOkgaw8kUq7W1cbO8xHi6euMsKl679
//w3pDnLB5Lf2lcInj/g19JU2zQ+Qf+bWdh82sfVbS0WJe1VY6geTGQKoewcLdbEXDrb0vUMJ8if
BWy6VkLa35goatd7xcduHzzRBv2357P69kAg6QO4yLC3cPJJfNoxvpy04tbBShNgF19XCnaD6WXN
q4KYLwW884DHsOYNpHZnRhN/hTVudTx7Mfs088V818sFoNIXcAxVYG0i1iLLWpE4l3bgb12p5Cjf
9Rdnx2aW103HcNzfLpZtCgsqszJblW1lX/aB28SGF+Zikv1lY5ZIe6UwvGjC2sTE/6s9os+4d8vz
kSHlhVk8mSiLhZWAaViSkJOkfej8qL6+v+niTkU52gFckcDaU02L6iqUi5vf7wMqcNiUSIfBhSzP
57kiUGux65NfStyGOm7eUXvvG60Goth12wJ/KimWuH6QcJLfnHneRMhIjaPCTbwCqE9hZhAzP1E7
PSxjWxYeyu8LAI5Lvibl56ykdHHGmJ9n4WAdMhtTAC1QSwrTO6iqaxoj9b3Fg0gTRUvGiUwwzEVS
wBt0ByqBZr5CeM5pr0VzHsRCZI3gvoKz3PJGSkktfgt1+MTlt+Ggqn7E0pYUNq7oYEcI5eUtdgma
35KhOjp/ntMa1+CpdGPvIKYYFvnVT9uGqNOGPIt/7c+9jLZtmPim+sbFclqQViCadK9CPOaWNf5B
2qSQAifOwr64VjpxaJ+ydYRWAvYUJfGsRSqqe0Q0OlwnvO47hJGwRXggtkUfJ+cD2q1cXrVFPjyJ
cQ5N9AXnSDaB07FyeK7vxdQXdqO9BLjciHgvK3lHb4hU45k6rIbW24WOmzjYtzpwZmkbs8xLnVit
ZQFNG4zCB1Wdqf7xzTo6o40GmLyqV2hJkja5JhD3h/RevZAYYayUwFi0ql/RsHn6KT/orkxO6jgV
OMMxlQBnPoSIyCAUiOu5dPpX8jPvOIcaNTVueEqZtgRWewnLjZ91ILIL8Hxt0XN6+KTq0Or7D8l3
76qEgljY3rOPXIIUnMx5l4Kuq+zfjLtj20ZdsaYWnHa5MSDcBrAVbV0P9XszJfx8EjjHvKfj2e7Y
XUmKDMJ5O0S7hMXvg2SdgjGoy9L3+zj4vfHMIszQwtPsmWOmhPFm2LNA/dfCA/fa+Vdj2qYm6By8
BooO2c7ab2pcgbZACSCL0W0XRVP2FTJFmtXez2kbrbZ0RKNkODlHQstm/HOQgemoeqH/YWfO2e7d
EkAlrT/mj5m17WsmwTwRUqz6owKioFuIvr0W1PXcgxuGvavo+FJMA4FULMHRt5WXSIB5j84IhfaN
fJKD786b2nqIfYTUQQSO89zIfqvEU8ssD7D7vl3WJWqXcvYDGu/iHdgaSZD3GUezYw+Ha61Ayf5h
VWQ+dymudAlkJGz+IVBB+l6gq5e8WfGd1Lr0yK5DJShK709MW+f0c9WUkwktFR/FkWxjlPNE6BdE
oRbIVVr7OOhwriLyGWyMX1vKy1VvcyJJl0epAazGj186DgkjFNLxpmkiK06dLQdj/1TcXNsgUBKJ
ZB2uRugKDqohIHS2oGdigNWUCoVOwOWDf1TfrSkRtK9E8dNRKKvNgMaRRA1rtLsBBwcgn8pyG6I6
TNlWGFO4xodf/BNVPSkbArXFs4wiBmWn/XhcE6F4foFgFtkCR0c7hJZj835edKoNhA2+FI7QiY2T
9VU6r6+qD4nTNASThrOXnzcqRluw74xho2AoLsKUdzmd/VtBLSXDXdvgi3EZL8wMxx8PKvRVFaHW
lZIvv2/YclraSlVW1UdWoajG2q5wZlbTRo5CUfmZ2FFywonUGOJ8xmKj6uEenYAkb+uPoLrTXyRu
kyQ5upZbYr8quyTjOj/qahdXr91f74zy0KGFcFP1YaVLr1+C6hQGHlxcqhDvfs1sT8BDL1PAoHgX
Hz7MsoC81l3soJNv1rPhxaXIdbgk+mwT7z/iKSmeOVWVzDUBesE/mR7JOi4TbK2Zid3cJcMliXbY
iEy9+dDvNra5FAZSgYXK7Zt6mfFiybeOk1rrZaX9+8gEQ9opcZLl6slMwJ/UuJy+hQ5n5RR4X5oy
N9jQWTE0clo5N5Eea5gvWjKgoKHwxmJtTKmg/IUkvQl3iU/2zu6pR8Rkn5qAIkLR+81hkUGNCECf
YE+6aI06lwC/3+aN6+pHtX+WUM9K/L+HmhitIE7dro+QCZRcyBLwCb7EuEv/APq61OBhQ+XgT816
pVpnP0QKcA0aFVfJbxbAIPvnW+qSeKWIFtZKdwKEebsGu19bAIxyA9JfmuQsXUJkkepX8f2VIcUe
8u7noXUErrZuWGNZM4TwMZyUJUKgwVcAYXvbPOWmFcQwC0FNK1gHiQ+Vu5Og+u22dwkohLAl5/Bw
3MnaeFbkkV+c+3uJwdVceSJzogxaMWX5rHaXyNVWWGw4eGmiPMq58IStJoYWPE343Q3U9prYTFZ2
AlxdL7sptFNm8VBURCC7HJQEFoqnv27bScyaa3cQPYUMLhQXYAN+HGO0JZXIXgNHCOEpGN8LxPIS
33vWVM/r9IG5m5azFZL4CeMoLx4j5u97e/tSGwCJpOcLXVzIwCuU13O+XiPa1MQrQs7+ovMlWet4
jF/IBFtBmASlr5THLWUAuCze6QF0iSXdDmQoyvztFjeRFDVVhaoxpFKaCAYGITrl3KJCcYoPtAkp
1m+86w83DpiUHFh9SbwphQwrKJkKFCwUYFy744FcfuPdsp2RfdzA91NJWITvqZ/8lD5xpDG6IA8X
oobozVuE/XLJz2m7wlfc9smOjtNfOkspe7UqahWhJflZYi4MZP/bzetIIEc8BeJ8coKeu5jZy+MW
tGUmpuFZh0+YxrOgucWAWuinmfMnKIM1YV1OJMHO6WTcDSOjBw2xaCRDoHocniFN96aWQhSawFh2
nkgNc42TsEl2ScElf55OLJUmehE9SYsTErNV0TT7QyuGeFs+rNWo5Hh80uDmi1CaVbArmh7MX+Jb
2jFyoiPEH7oASAIKlzSbtbKokR7p4sgVADZ/ZoEYwm3VawSal2p0hLJdeJt2szOW8sBj0Tnp0101
tlxzh1T8jhJ0VfaMk/aejmcm5uWKCYKbW4SFLstGWa8xzdNPrpBBVcjNqPs8s3r/tRZhkjnsb87I
iBIfCnmaYei7FoESqfrGgtpN/3dPr+di7yVaPRJKsPhZNoYeYhz4DWcbuchk6D1rUZeubv9c7ZdA
9Ra86TvXqUq8t/3C6TybwOGh7nDnE+IzH4lWyVPqJH5AvRu1MVgGmtcTEWCkN5SQPb0Heuh9y3gQ
1hqA4H+TmZlOng0duuwK1UY6WYtjaQ+XH712QrwnxQNf2Jv6wv/jIMRYjMdFgsr9oXOsByRHHHNH
Yne8TBLp907EUyBTIW9WBvCVnHM3nEyf9a60sks+1eQ8cWtVaXxrAz22LkLYll2lYjvnDE/gvvYd
2lRZtkoaIHy9av78AJm83A3hshywYBDa4SxoAxWue2d6ODvyVM/JERzZCAcik9+77uVcj0xwuznx
g6vbkDr4NyQEsuKzppEe3cIyOSVBx7sMKHIWKOck4xcXnToIN3Wd5xnqd/lM58jZxLGsuu5RZu7X
RXJgcm9gDyUDZD9OlEg4cyrJEyVpsmONzddiXAqlY9pjxjF+ctR95RF61ZsggagauDhRe0mkjML0
Xn3VIIiFYzhf+YWZNbqk1bEnx4Iy8FB+MqTZHiT7gj/acCUqdh0K6jqoJYw0TGm6nXE6v6Zx95Wc
sz7dvembJDz9qYf9TvNQnoxD6wROHFb/79kqV1I75sCrfMfcOD9/Wd296iLKE/NX1Vjjb/xIH0QA
uw6a0sgtjJqvmBCG3Y3kMoXJJDJE3XBK8wTRumAlpVxgN6KW9t05HA0ohQQ01HIxGn+wmD1TQOP1
q0nflZh7Lq1bznOQXaMZAXzvTqehFaXZMGhs6a6wn7hp9DXU+S6py4IlADhbJ+PyTkoDW5hAv4fc
sTisnLJYw7lgN/7rrkcV/SlGCrK6+XPVaImDMM5o7SyFs/UO1r+e2npapzTWvLCoJMtDP8j11UcG
xF9mpFgxrT3rLOz6ywi1uyfb7XLtFb6g4wM4ZPmMaKPCovHtKX9Hq8IRSYME3c+daLaKXSxE+4Oo
6UHjLp0vyT70SAahvAB/IwwQ1djrwwr2gSlK6aMpZ5eFXpIMmcKoGTya3LidVKHFYtHLTaBZDU9F
PkaFJsnE+6XxPDIZeFF46YjK2aq//7t2v5hCeE9/FC40GNOfGX/DmgHej8D/4WEGkF1+1ACP3HDq
8Li7WBF53a/dNQUcO1tsi28C0i+YPOrLuZfmMJUb7ylfZ7dLJYtPpB50q12pPqfxNORh/g9NkOhZ
At9LygaCzxhgqFAlC1plBW4sJc3RKnW1hbpecwrGRL43SoR1IHPdCpYThLaTliA8k46oschItWgy
7vCbjX+2cP8iKyIfGQx2SRDt2YutVgOHDNrv1gvwnRGRGJiaUzLuPLzueGx8cCxQ2rMaBRjdXf5v
jZJganUzJ2q5RR1Sidr0mICCOVBB51VsqehUR2o8o2rBrbze2ZSzR9pigGcr82OII/CoWj65e4JA
qKun9vMPMjLYpRiraTtNL/eKqe/FmteI9JCNs3VFXqD9wBkwy8HzFRl7RyN9VtymspvixeX+AgYc
QrHbvzxdaCQ2QUWCyYjItb6LMQh8cnrgfZr0rlbB9IewLRLSBuo8lgP+OYWIT7rLyllQsg51AIEY
vGFT8uXVyPSbub8j+QMj/9NssPn+GRynnuLqdv8RLEXv/igC0CGAdMDXjlbg30Hy1h3nO7XZr21t
78CLUDAxp97Wrn7sZvxEi0q8sdv27axADaOYH+Yb/YNR/LGLsbQjOnGV/rNbn4mAc/TVhUcbtyk1
2IG500lleTFaV6A5Y4oqwn/UrpoR7X/Vt+RitldzdKMKSPzrTsFSFlw9wEF6+BEjD4VcxNj1hHkc
TUvN+Wk4aEqAdVGDq4iSWDnSAKvRKWgcaoQIxh0ayuiuMUoeyNQ6zr3xt1TAZagaaYGrjzuTacih
Y5njhfEFk0c37M9RbuLktJR9tPdzU/OQFE7kkyJVXCY/W7NVyk361Pt4o+K5XWSY1NYTzXzJnxF0
tj6oe94XGvmOfDpPOtBMj0joToLUfw/vTOUm7tDcyK/I2NKLyCxpsh3HAOemDhHl3wtIZ+csK4zi
dwheP6hN3qsUmwnskw2rLXiQ1g3J7Z3ZNhrv/XjGkOcxwuNl2NQ2giQo+Nstax+Hm6ph17AM5AHS
gj1yFwx5kfMOYrij9asSl2OhrFKmMhnVncD+QtqVnlYGVSrzVcRSBwlYrA6aAXoPBX+0DDTeG1ec
SqekOdj4Y5bjnQ5JRk/HMklx9b9CpzNG6+6Y+QPpkpFlYe2OHj9g0tiUxsFo1RPmab42HXH0Jwy7
fZts4njWajeyCsF9PMJgKfiI9ms5t6p5qT9CvSTS5sR41JC5UAujbfTYKPLCvt8cYNttenDZBV4E
rFPbPxGamMQygTdxGOSTx+wJGmJ/Netru2mKCDsq2hDB8K9rq7iAQHvx3F2JUecMe9NeRMBUZ7ar
3Dwcv1efvdUuNWIMcsnVkHU+QOcHue4FqAgw4nhhIMKjI+wlPJ3S/fHTGfegksG+V9qky6A6TKlk
llgfhieVZMjHppIgaTTRdM+n5oBg2A8DHAZzUgQue1LDHVDLTotVD1wXlh/N4JbA2menhSO1dVzP
rSR+uqwJUjB2otDUPDFes00oZisMTprsLF7lddWY4n1IhrvEu8XSSYJKcBqZDwYNW/SCDcIyJVuq
hHka7DjXo1/5VcXbPQW3LkFu2OXSd4EuuRlrJFyp+RyYnJnEwlyPcvIZk/qPrFpF8+dadAVq2rd0
9kUpQgq9OiJGywD60n+zIgh71RH7YTuQR28C6+vT7gtCXqw9rqVNZczpXBhQoFzFw1zQ4ecxGzRh
nEEr0T62MzwVpnMsLhtnNulS+JeruTDogw9dlKJOSG7NfEPu9RJH/BNAJibKoCmhs7xURXk5KDHl
QefKMgSP6TwuNhL6YvZzuhUz0FqzJgdez+W/9DUzPGmWHCm6tGSnRG0IkeQxDqdDQaHskph+Hzcq
4cqU7cY8lL1iAFQbFfh6YA0Y+2K6vvKQYxMIe+Fg97RfojeKL2eRjJT39aTSBPgktPwdnBkpoE/l
e5CXOocsiXYYYQejb3UorB11eUZ1Jt/DP1CBbAicu7DWs2umfdxQ15BZurC+5bNVoK6hvnPqdhNR
f7R780/+F2aPuBMZmfRxV/jPTZah2/XYb/rpWqTBbM9X0/tGt4mnXOjD6hd1YOpbAVIs9CDh2uV9
TYdehgjDYHlGk86e0E3lDpGT66SxsjnTfsNejpXT2TT3LRcczD8ADwt82PgeVExPf0gnz8i/DsCB
I2x8O9Ss5KBKPWCSDjAPcPSEsjj17wEWi1dHwwZHLtAeVPBZ3bK28Wy0MtsQTibOY1jky3ADWBzG
QNtrIkoIvWCX4dU9y9/X7e3KWYoR3fEPH91YANDhPd2vmDdgxx/9T0fM3Bee7f9m/XbBs40bW1La
Mge+kn1dgB8nL98ohwVkI8wIgF1ND5C7zmTHGsmT3H6y1OKnlws0bK/+e8fyBp5FkAGBZmuGak3T
zal6ngB8b+KG9s84M4F3Ah8YgIYRFzX66aFYhz/2P91GA6Izpi1OdBhBs0rhneODuUtxblLcWuwj
6et3dLM5/xLIktf00MPTN6ruMaVm//V0+BfsHMktYJugWPXAy3BuC+vCbVxLbGCpQhpYJ3dj+dwy
o/yMLl65gItNmaOXEqz4gO8KCo079SZdrTV3OSiMKbhy5V1pbZ2eU/cvcir85wahrgUeukpUXEYA
sRJ5sEltjCRi0ySdaU9GRMu9wp82rRV+fK4kDu/PggdtC3Sog20dOUZXMMjrjFtOJE6q4v+eei1K
/J/Vq0XbHkt416vygm2D9gjpum7JsnlYYlU+Dia4AqvvOrLAOUyFYKuJbbK1fyPJ9MwHz7Whs3tu
OXYs49PRSOTbmCDYkk4CbikqtnvnXI6M5Ve2Gi1rmvPsUIs+AWPSh76MMOjjXOf2QyQS6JjzfspP
kt0+g2IB03zFqih/ZBCg2bwG06w2cCQ47ioTIoddeJIWz7vspJ8bjWe50SKnTO7bGJLA09DSLBY6
aTPT+BGGBSn/WZ9P/CwHsNxnFKrzQU+Va832y6DW4X6YnxLZqIMuo3NWCZ6HGplRwVyTpGlobic2
XzshjEzxGBcSU5yFV0fOxuSCZE1rME+mk5PHKGD4VcAwIpxZZQQcaktWmNA8O+OeBE7hRRf/Y8W3
f1YtnC80T6Ffzmfq688aNDrhMGqF4MfZougRpPWERjA7zRUSIPZnxJxpF4vyXFVJ6rgH2f3XbR5A
Pf4dJK1bYN3jkGonmHC0UWZzNDfKysXVklnw7C9lcQoLSYFLXladbmNo/VwXFvkdAiUFlZ6zuo91
GRItUBI0+lp/qDYdmwYexDVJ4C0dTep+k/6K0ydYI2JWDsTBhMtRYGXbRfcHXbggHNunpINqOq7d
GbWpeN5y8Y94Cp8Kb6oeSltbXqI1FPj9h+U1e8IUSt2wRG/6QjeY/9SWkED5X1Oh5uvhd1BEvIth
ZReCP1F1PW0khyMnI57jOAG4yq9L9TUrDkfoY/lnd8kAenFr4U/j3ZoYlaWq3T/hSyBJDuXAmlOW
1uq6awDMGK9xbqQLURuJyraDpwSDy1eAS4GBfVBgWo8t83UBkdH5uUI7S1C9hxitE8pYi1UZoE4N
nNSiYn5DIZYaRxpwKXbZCjJEbVLHADMCwhVsYHp/SKp5fM9dRQmDIU0GurvRKgl2yCnrCKRFGg/d
41w+Niy0r6+7WwECE0PvPRRrFE9V/pJOPTSzS4cisR2NG3Yyu6C6ue5pbN1fW9KIhgDBzdlDPm/q
GPhN63wKPME5l5si7wSRDKRwKgwvWhjb95whFCUptRxT1JOoOJQpyw5GwAC32oEdGKw9gIGlJtCL
PkfcDiNgVTUqWL8/d/KM0M36tWxcU4mWAcjQVxb837aX7JMpvWgzsC2dDscFiFKxcsOQZG6btrfe
M5oVzCs789NzXZAMTr087gung1IxxxjXrcop1gRPXHzI+yGh4Ax/9hH3rRlorEkY91e1V5mt5x/v
5/dAEFrlsHZUr4RMviBNa75quC/1pRh23mimCe4eZsfY/BPdpndguQOzo1gk8IH+T4q26zoeiY1d
Yqki08NwuTgOYqwwzK7xFnAFjsyON1zR9gLQRZEMEsaDJNZhaOiQ6vhsHqVpAvrtbVX48Rue4q8n
4wJRKTHD6sfXLrRlFhDWDJyKPpakKMKjpIcZ+BBMrNl/GLHoaiuIsimcDNGt6rC09wrE9dhSF8JP
zslGWAqBeICd9QJBgqBOzsD9sKEKmB7ilA/j2DdveDLQdePo0PLl5xZ1M2PBfwS8FzZhduC8UBk6
QIhClEm2m8ncw4a56F4eE39dvsJS2HinUHfNZoN56PsS9GNdlQfc0P+CqKw/CZVHt0esMJ0C5qlU
It8kJYo+VEBYe2ihBrYfmblTyYMWzWsRAm6J82VMVcbRYesSPJACy7danG5LNwLKyBJlrIU9YWnl
2FvV7dkX1E6n4e3I5/wzIYNTiOu4XtSFomXcp9xDmZS5JUOCQn86xAv8BGjoJ8o8d9D72hhR2Gb2
U3gS5wpTk5aHLd3mHJ/QLr55g5svC9b5IebPrrZcZAe71gXQ+gIMwV3m3ykNS4So1EOeYI2V6Ats
R92p9kn/HtRx4ovImWHAxLSDaaD38hON3DmcU7w6qvfVhEZtlc796PT2HxBAlUQ46MMR5VdzPtBQ
3S/xnp5f7sQoLlefaEkddV15BuH2g1yP/joXbliQ0SBmYsyMw8aBI/OHfj/2SnMvcKp1TwR/H1Gw
jAQ5VhQA72uallKgeA4MmlLEkLBm6ACPdUWuOOFOQjuekL+gakI8GmYF+jdNr6CEIZh5qHP5rx7d
qsQKeP8Jh4sg1B6aru5VKE8lO5AdYiGK4oWW2R3eFaus+vLn99jW9Tx7lgnNmuu1cXXcGARMOnhV
2Qn8OgsiGWvhrNMaE12Jav81I9cBY4ZZPfO2mCEGaGuAxUdPGxAP0D6R9/XwIeJ1/Z34eeQVeeXH
hLVxRxHjQwK6FkT3PpL0lqw5krcuxU/n9OVqwO4AqDqCNB9tFzqJg0Gvz6jwLOgYL9AuAZMNSbAj
IWT/TvHTR2MiF8L3X8Lnce4VLtxeYKSXdyWyuZwfNvNyR86s+WVSZBymiKBFOEtagCALGNSaCr2a
XUZwBHIDqTME01zNeU2PXZUMmxmhAZ/bZs5QtjCO7UPd1U34PI7qVp6P4eLuBscsXt9gfEKccN7y
zW+9I20x26W29JMjWNoam6FfpJ0gJwPJpNzBxNxc6QYohAm78S6PSPqmL0k/kKR06xLS3vq7efPu
xDLnkyRuV/1DkdTMNILnSHn/K+jnr0BBADa9COGDsN8pyG9xrqC9EYy4o40mil2qoMRmW/c/CgaT
gjUnFm5VanOxzZt5SLSpaGbKu0xYuP8+sSP5jzvtroPVEOiP9nkQK2Vkph6qoGYQs0fc7fONnQPE
1tS2il8ZB7AaUNFRccGzneRICA9ivXMvAc0uO71gTpDz1DrTybYeTg1dv7YwBfNUWlCa5cyuvCtM
eWh52eRLIXjtk4fmEs8nuPj+eU6o9hWa/XHkqbkxxwXJut5g5SlTmoZMuItYu1hDh8z/8khgSeOQ
GRrMdtVeTn6a7BT9IGIM6iAtfuclyz2pl1gVzNpeUgvVuO62YoqsrOwVcRgpjDENX8hMoqtml+Ym
6+Wa9h3xZpJlF6I9aGrMbWhciuLoXtvxknRwziDbsPMmddjRCBCpJPimyphMqtZLuE0f1LWjWWZ7
mmBkRi+QdX3TlYUGWjYDYlEMaKhmdTvbt/0391afE1kdNFBwxc0OLi1W7Rf7Dc/r1MMknNzLcHuj
BvVYs4I/8+s8UAvc2uXqbYqZnxUafR53uidn9q+aYtkfg4qjUr4igWy4J2SujtowmwhFzp10eool
fBGxsFd07E+4BwQmJKWaP1qj2TMpmbQArx8nkyRNwE7bx4TFOqfyZUd1M7a6P4wThrPEXVJwAB3d
oQ6tTzqv8UaqBDY2HF19ZUKtuGavfSbIfn23qEC7cjKQORu8vMH1LlzleL0z4dbGPUN8tlCbPKU9
PeJ0W/SYqPGqSbAE5Xm02VhPOtLCPWA421bWgTL5CUNVrjW60Njjdq1NRzCFNyVZDBC27lTiDbbs
c82VDowRrVTIWBsXEDuKyoBeWMnc2dwVHwlf3bQgmKxkQxw/sk3Sj5XL/mcdg6e1pLPzF0ksjmtg
SGqPmP0oLddp3B56N5K7tHDW6jGxP9rsNwG1H/7S9gOkylnGrUy9wBxZlM5OA3DfMhOa1eGYzzNc
kobEa1owkfp0Kd8y2iTXO/9yaV2hsGXq7XkajGuwlUY9n1993bhlghaeD3hrYjwX8bsV0FxEHTLs
EXyK5TUERpuUZOEeenikXfEDGu1Y9tS39B3hJn2dbqgA+BjMmxUzNgPJC7iIltqdhsEWubKOQ0XT
WiKJaWZP7Mr5hEJLnlG7MrN+HsI+yrlLxjiR/vD8MovEcNNHLds3c9mpxYlB0wHWHNRhVzFCA2Zl
pzGjXtTNSJ9Bv3luqUfEUlwk4f90JV0z/uzJVXkATNuR4NtHJhpSvrvDShENlAUAx7ue1Is4L0TQ
25z02o8m5/LRJAkkbZw84kY08LSQ+CG8syiJ9Q5YZNcmZprcUgtUDdnyBpnzRnZCn6UQ9UMvq47a
78nOcMa41UlZIYt1O/Zdq91bxy3+mwG/za0jDNzHhxRVyNr6I9bAGmsZfsjXayqDM830ABVh/PjS
1crvZ3/vhI+K5wy//zX6ukxNoaw97Em/E4jTf8hj1g3gfFcpp0wMOLnmsgAhlCLSH0Kh/moeFI+Q
Eh6BWnn/CwyQl2MbQYts6RnXaXiw75OOkF9QxlO3hNW/XQz6qIozAZcWQPZYhoWpDXFRod+4hRIN
3VX+bitAPYj6M3Tak5w9CBUmPDi38gOjrETLivJDo8yKzQi7XMISzqlFCHiIJlBFSuM/kqGPwJBR
ELDwoGvwR+aEwReQHYLw8fTVxgSwH/Gj3zjF+DcvUTTtv+abLYJ22aCrq6q5VpG/9C/3gGnc7wn7
ck/RnmZ5UJfm69JurTDtfo5dWuZflDCZFQGkccBxicoFjqHoeABw0dOD8xoYC50J7RNyRnU+38XL
JDWeTzSbtN6Bt+QE3AQ1sw+CIQB6hardUZwCSU6+gk8TLgvOC/dXb+7fCWYjBBPTylrs7nLlgIu8
9WkMUxssMyQRUpDZFJ6MSwqJmRbEFhL3x+huDhynPUcAwyfW+GxKLBo63RWJDvzGs3y3TpPrTq04
ncFfc9ayiDR9VV3ZrGQwCLoOFAxKerkRXBhxir6U4rtPhpGyspwByZTCLT+iIEytCpTy3V5Vm3yu
dj0ypaaInsoEoUFYarMY+P3UJ8i98yZzFuQMK7qKPncIsHqDB23QKo/so/jJf1/TZ1VL6Zl3kE/5
SXo9mxF3yS9bbNkwOLNlsiNYTsK3giKVcJpnOWPpKMlrCuLQMfmg2ChDwy2oe/vYADwFbdscA/F3
TORgAoABcRIgBI0EQv0BlUzkVmdZ230NhfSZ8WmBIDd+Sc4v93CcGvTVGZl2y3Js/2XPpnb8prBH
bWcEFO3tl0cK3DgTY2BZn7A+akCqNAGhdXMibFwjadkpxza2H5Puo0SodeBa72LOQHuBrh/T0HQh
DYmGPr7l1IvxEZtnku3uBG5+K3u6Giu6geYy6zF+LjIzzybCQLyLQzSi7RvoaPIILFFmXI+4qne1
4B0rLifRNR2Oit4b6UG78vfGKEWVHMEdtNnUxEAqjuvEHxIDtifjv4TG0h6kbmUlJ1u2nweNZDw2
K6KJxpsInm83YWRocmLafPHL15C40BWuXxiNcPT7wShRygkFNOCUWlo5UsjOYklE2OwDFpXFLxDH
rwUIUeQlS6WllJ3c8tSFgP1wBR4cjI5zZcxbj1sS60rm06CMwJi1KU7oIPQGRb1/V+tLxES8GsRR
DU0hK94zV4js0D7pCtzWPk0erkRF1AnlP7w3wdJ3GzYtQyM1zX4kF4rMuuDnS4calBJyHQj8wgMV
1tSTZ1wYjAcuhF9MPbX/gVAFzhhYtNqMV2FaEMGciYIejICz0ApoDM8YYOB0HbtawsvLH6044EwP
e0Pu8mGhKBJaOiuzqpXBRbQCAgyUSri5bg9tvPryaKkJ7O+T5IIhkWNcfHWBXx7qlFpgNmn/i46X
vy3+9qfPMpEd6IloNmFIg0lZC3R9Kq0CwZEfkX7OmfvMG7nQ1QPgUnXGDwF/7iyKvjyGR/YOKEuy
ETh4LkP2p9Z+A6f7SYsZDxvxB5EOjlD7rRgTwk5TRrDfzjrMEXJKOWByo1lWMPf5HOXBBqzB8230
eWEtwyivITxfKl3NuBuQj5kHCEisok/uTgANqUxtITd/RI9X0ME1chiNGp5OB880C8Tw+oo+USU0
+FL5bHj9606KBuHVHwU660r45Gm/5Tfa1By91qZaRvUbv6B2ar1feaej6JBy/m86ZCVgXgoCaOik
MY0EBEC+mHZYSBeAoim8KJoUuF4Ao5oJyoUulQNBV2NL+tdWfsbbABJXfmnnoNvhkBfa6v1uQHsq
ySp/ATVM3H07wdAtWO4QjPCF4e3DcGHMr4aNH9O17tSYm/dlGysZr81SR/bzm+VXVcPCNA7W/7pR
2wmzzD5rpZZU2SxuTEFBmA1NSbyO32LiIe7IXGUqxCECL8+yhXZXigQV8X8MXVc+4A6b0DJGnl6k
1c0Otjrvfkmwby6cIOLMFzzcWUziRRMy6vDNOqzlCieeH5l522bSLTo7Dv/cvufcTBTtyS5hXbq9
oa4nuHzQKI2+PnfKSGDg7FK4i3diFAkqQm+6GbqAYWaeFa1/UPDoabQckKKSt93sBWLyLk21tDiU
AFBWO9pumzaLy8WAkInMlagPwHTNimGlv6pXLfdMheRrRUfouymOVcF0Qm8iOH6gWwubHjYjWyS/
qn543Hf31inSfygaVRYeYWhxe0XFNMEWLPbyCkD+o+99e+MsxXPf07f3Xk9apN9rRkjIHnDQ0dv1
fasmGMK2x7/mgtN8prIgKIpSMSpCus3eEEcMBoI314lDls1xXokuumpBDND2PgFCv0iKlTFY460r
09iwzZX7s9f8bkdlsSZ/Jst5T3k+ERJn0HoiATFf51zOmIihnsaXIZGZ1N8R5aifYZ2DIT3H17ei
6L1oCdCqnsO6FiQDS+sIuA7mEy0sWhFzcrZiivjGEJOz/9lh77H41y1fQ4NYhMj5jVoz+qL9zENa
3g7MXd1LuRwUjgqzVt6xeXfnZbDIzkHFgPPaB0udXvgKi8G/fGcXLChTQujsH5K1qJ91ZH5XbW8h
EDP32nx+azOyETOaAvejnKACGnUrVpba7ALW+FIQNkyUtJAZOmJRk3hvxGyo3CxSQUCM309CpfdO
ZWU25yS21YeHyRA/Crn3WfMmHMrNIJmlY8KoIQybSK2DfqNY1aZpPS/MYlZapQ5L3uNHqoX/ZE6o
mWXsIanImLvXBqBqIWZQ9EBKuM1LHugCDrfvEr8/L5pARSBCX4Uj6w84RoHvORdc7MqtdJ/oP5ws
vth7Xb0DA/LPQNLwzXXqi3EqvCafQ66abIjCsg1/Qj2EtHNAuOOvhZmzpW7MDywyztb2R5NRWOhB
50VRJx9xJtrrn6/g98tQyxfdAgdJaA1zQ+gteEdajFTeoQsSXgcMuiv02xucsoVgni8RWGqLD2/W
b2laMEPNJsKWEX5QCBbRJm9IOeyKjtaFIiS0awUhrl/73gp1/F56QGBMab9LDcPirfyzvFNIKS1s
qZNLPaOKhZmuW2xqR4ek2rYGI1tEwCy+U17Z/V4FAHNv3qa2hJQiRJ4SYOZoC41aK8TS05XxuAa7
K8Wqy4QRze4dhP/O9WNdRp1yHvIaVjDoUxLit0vbfsh/T8Srxe7JKTkskmhNLA1B5kmcuBk5RXZt
qMHtdXpm3AglI6/pDjYFVUUq99Ptxk9HTOut7P0EeUN1duT3Q1VcDmTiwbNnGbT8tWYuq/b7QnKi
DER8QAD8DrMSjI7j5QrJnsMVcv9z/1a47qgxIDSGS2d05XCTL3lKf9QWHszDXER5LJRBpkW3Dh91
JW46MFJGA4bg7QmQOMA7mWNHNwndrZo8uoPDutr2jkDxESeTM82pQPMlZrxTzJ/zKQv5+ZqEMbu6
LwqggliwpGqd4kBT7wAO2xFJQuVq7X1CTPHH+JNrDwIV97PABf8tFjI+4dNTUQOnLipMylWl3lK2
DhoN55E79XdIAruvWzX9LemhE0kghOWVC1CtA7Q6pJ32/D5+mEn7cim5rjjEOQ3Nl7ehlIDullyE
5BQgtqXBTPYb/o3ADrYRENiEcfFm4yEzZ1pbb3HNQ6wwemzaZ/r71dno/BAvPRZyOJKgocWYi4Wc
9zZaLbRp/Tn+AHI3i3ttjD6WPD93vZBM+WL0gnBVLQqJQDZIKlPppPhD8ENjk1N66cmUBmbeQcEC
WJYjtoyJDqpfbJN5MTb7KfhLo8W7XDKjb7t/QEsPPz7J8UvMQm5MT/vmmwh9L3VzPu7Gs3RudGoy
tPzOYb7rQ8lSOwcZXx1F4Tq7BYJ75P7rjT69EmYFHee2cEeSXaoNYrKay1x/pkVnc82hGJVlNYpf
VEpdPkMOJk/bhUpKrbx9UBTafKXKMxzFR4LSsHGD79PAQfwk4gUP4ca7yUdi5455OhfWvq7DFQ4L
dCl9RFO7ZasTHQplbtKwHzayJjpkdlD3FHy3E28KWGYqeQglRxdZ0Jl+AMdvDGqnzTo+dkg3GL8X
beSOxlOjPRRW+dvcuw6jrHULYvM8IUXqJlVt0qG2tohc2Nd93OkXUAvJAaoqX8lrNMwOTb3j96CS
R1Fs4/PfCHDns4w7nrNtV7QwBN4cAC3+dIuEbsj9oPUuagIPJr5fxYKFXBs2c3MfKTl+5uxhWVKe
m/zYaAc+YQLzHtjAvkHsmIqIRvJPSrU3HFNgoD9hSS+PTt4LQurJZug/UPfvwC+AkxZk8WVYa7Pu
FfSThgNKbT/Li79jpic49mJ3N0KfWSkO73lPgjndqSPSZjxp/7qNj/2eyR/SDP91513Jk7bdr+wk
tfSLuosOYoZnzkSsKP6anjavuCPRTTYAJ21xgobHP90s+X3wkGicDIB5MehwYs7KJS5lPLCkNga7
fE5WHIIJiJJ3idt5IYkIM9AM5NBAcA97QpP/PU9WW8IKsKAerXzH6FU3H4g/ITkS87dZXTZcdoI1
N2gcfe9oYbvAywC3fcJf/MxyiSsDusGVPiOAH7KUVqVaVHHaDWOTJy+gSVgW2QkjNn1qLITKFCqL
Qrr60FzSfzNH3Z5Bg72qDTFx8a139w4qrgTZYtVdfEYi/aiA2nfCs5jgEE1NDkF7LJxlE4dAk9Xf
BP0p1yqLOSW5rPywTlKE3gXsReTw1X75wPj6/yoAZVU28M7VfPfhcqQ1VLKvfzkaPTJijNEiIQFR
1aN9M7G84v7neEz/gatqvT13Y7aO5M/CunIOz58p4Wlk6JhILJ1MdHhO2WD0AkmRRWEcvaUG9H50
N3Ddk0zM34ogIOmv+9KUXAMLi/af31bYqayBdZBktPaV6LLCG8+/SE5/VdtuWY2cW2DFetimsR+P
N8iUdq6vJ1hJgQ6roLOAL9Ncax/tmYIrzuF28C/J+Qf9XewLFfpMg/OhZdSNij/60GkJlaevwnkl
fggLrvRIHADb5zVC1qccCVgzRmIbo5vKV/Sc1Ci3bAVXo8OiioL+z1khNHjP1Bq9UEdEaW6WBzYY
75WSKfIA9tptM9kC7EvpRKnxbISbpbL58BhunLlGSd2DvS2W6cB+UV8LsDWcEyTc68ZEgTb5LbQV
WLy6v8+aTPDMDbCmHjw4sAryQR0T3xfghTGCIq+DOeQhFDablka9TMZMzlQJzp3xAswnfMtU6n9r
XVZdUFAap5YCB8pZ3f6SyL8SIc9GMy2bhd2QnHYlnLvaFCeknQ8lnzH3+47wz0js85ZdPr6ZOEip
Y9OqTjekBQHQB7IDfBc9j+3zMN8/ZQpqq7Hx3vyDomHuiK1phrryVFij4BbRDmJloztYw6osva5J
jKsblw2aJJqfcMoGqqX1wqQO4dA9A84JuFCQa9C1KMfl6tyXkaBnrDa8AHYZhTrXQc/LFSke83fl
zS7TH7H9rB27WVNvMDyvYVX5Im/SpBlblbg1O/R+YMHebe3dK6oq9tyE5SvBsLCecDKEwku0gXpQ
KUXAXfNmJalei7iijSDiYxCqhT6WUtc5yBNWrWdVAjVfyWWFg8AM6SmgmhMg0BXZK6zsVDdUBJdz
Z/hFsQPubdu9na2k8RpFwwu/b42sKrs/0/Kk9BiKvVuTIRTptMUVfQv27rZGi7yFXYGEt4MtzEuV
LNA/9O2PxzSh/mF3as1EkdNjCfuA1EVQiynG1LKljAjt1b1QvP3CsDdU59hP1XWGk+5UyQzpJ288
R5oZ2iRC3NTXBNn3MV64ptWEfnvVGgpjeEjfyds0VlQAOGffK+hDezkavC7idNtR8fJXVofGWjGI
ZN5aLFnHpOyKEwLR4PX5D8clR98qiPBvlDEdhhaHSapCqP+2r6imbdlrWTRQzaYieQrxSv7Qytrs
4Q9B6vhf9QhKXRlmECdNlycvPkkIgLeydUDB759KNRRrf2rmrSp9oolEqJv7RZSIRc3MlQcGe9OS
twaWPC1aygL1HAxmNuxbJ0YKhoEsSHaXdEQ7RPXVzFvXwmphfy4OtUqOLXVUPddljZl9aCh/hbTQ
jNMztd55CCeRfq32FSFOv9mrxCONl27hgAHB+oC0WmvsgY4rbPQBcd9nr5OtMxj7fbE0R280xWp4
S9at/Wya7TjwibVsm4NCyIA1b4tojj/lQSMd65etaggRVP0aTf7kAblWLeCGoTsvX46N8egf8Cg5
Q3T+6H3tv7aUudO830XKT0k+iKwMGLaCAVuCZEpfPQEVySYw36XDaLkRUTRnaR/YsMN1/3raw5GS
DfGeuLyCnQe5S1rWhGY35hALmAZBshQMl90kXMRmbhtFJSiddo5nrG8jbYY1Bg25O1Yu4XI7IBqf
2UrF86T0L47YDNlxgnfGC4bMqYMaPP/6ruKO9gzsPP3PnlVbi2hiSzk5BitP2WhWws+8AIhxpW29
JjUhuT/YwTI2acwhkGUnooOev+ELCVJgGrAAVGaswIOVEtnUO2g4NREmqZ+nd10yhJBvP/4Nn3Xx
0xZu0vgVwjbUMLFVgDlyzB4w9paKougnC3Ny9IyUjsbntaDQQtzsiVjm2tB87LgXOU6SK//OSCCy
PxfNCp7vyo+uEmfwZa3fODdCAgD2qTGw++KE4d60Avw1Ant59/ajZ/qMF3QQ0Wn7sBsWx4Aek4Nx
609w05XD3/PUz3c2687uPG42FFq5EqVwryv1ipVlaknxucg/ilgiB41mFWQh9rf0THwKwc5H4Xpg
Y2yJYvlJyID8ZfmSCswmC22b1tl5qF8IjM5gq8522C9XLsYJRojM8QdaDjE5QN0pd79qnx//6dBy
B6E8roU1TEElBXx5aZAJ3tAq5Dm6IsSdwTnI/7/wgJqidnlfXZmf2j17o5N7vBnWHrSOYh7Eoak+
EwDPqgPiHUObs6YrCMhRH9B8k07ByegmAutcA80srUvAUSQ6RkvTMrNUmgn3dhIEV1z7TtiE/NgC
xen1hOlmC4vKa4LQKE7reZigjooZzo9lzWQhkU51XZOjbvkYLWCN574UICWeryRBy4upPU7zhlgj
YqovkQSdchTwz1VhOPT0c4C6snKCozYjy5e0UoVTcsEs/R/GAzJOS6egc+nxRD71wiV7lIJs3COL
ld6QtYWKRLrHm2STf7OhVx17a+YmBTeMhJVCWXpqhm2B+j+oc5cIBpUc1yffGSG5hgXq3OEMtX79
pzbD2LH6iiRE/JuFHSN08T/RHnq+8fkKopPs3WufvEe4M2DaRnDqwfnqCIIsEFz2rpBYgOIkBvX/
dwuWsYqLY5tzTigWCKb5MdhIfLnf6mCBCqJoOPhWXfIfE0GzaQTyR6HZurfLtsoN7sfKhF+DWGAG
tKdf1lhHj6uSwoZvlTg9EYid8b/b6VajZB7+jM8cpHB50mhOTmDjSXa4VZUsRwkjHcZnhnIJHTda
j8ejXY9jgPkCzhtK2/3vCLejrYQM11E40QBsY4R4ABnPBHiMQ1Cvbo8kAwRcGYF+mVZXB+B4OC+7
f5PlkLwSWo6nILRRIwDjcnEI8Xrbo/ZpcKr6Np2TG59323I82IOxtzdPF6xqt4vlfpAd+KTRgBy3
F9DlzsO+wqdXiS4LGnlGRVNbldITeos1nkVZH53wZNXOR2z9V17koBrl4S6OQOqhlktn2v4F0eqb
tSCZT7ljJMNH7rBKTgR3TuJ0yLc/2vA/x0dZMgpxT1Qc+wEwKKJf1/laNGcjLwBYH2bVSccr7W2t
Ji2XisLfAvlO8YjKKaZtWdSbK6vGRLl0rTeWBHq8ENHmzmPmJGciHdUYc7kqWKwTGrJ7dh+DirQd
5sgIfekGHccHj4CBUg98Mish/v/ROw7JHmjbQxOJ3pcf/axq0AcUyQbGersnNy0MarJPB0tIppmT
UPKClI+QZav7OnJlZY5JvIiS/jBNpx/SaKVX+0OBsEl8/ypa4yTH7PmXZ87/AX1ejVyZVE4UwJZx
IwwvqP/8nr5KDnH8s4WbQNP4LEIvXNEvTKEzinchpSuSIL7fp1G67abkyarmcxWsnhcF403JrXU8
iIWubFPvOUhZqm/DITmxwhXbkGevq9SC1Ek3OB36A8D0oEG3x3Jjbf69jPzGUEbzPtdgZSvgTqq4
WBsju92Nx+y2AuYJVvoV0h0FCflnK2cqMlj+tDyZDrUJhr7oNR0F9SNTC/qnGg1ks1Y8EGBoElUH
wDThDMBlefF95q85aC8kJ50+0NBb4Fz+H9Q9UTQAQtpVgU9HDo7l4MpzEoBv8eL2wp819b5YKkI1
T8/e8OasLNjl7H2jF9lqKSkyuOdlsNjq/bCB0fFV7a+p1LW5kPAvILvGOwu86YdStyBr7f6noYab
5dWT9eWUMMDZAWAdGNjLY4gmThoElUUvGn71BxYqsm9ZOk9HPpwTPp7IbcWQA7st7oxENgd6ESP8
N3aFNcrmbJGbuozk+TCpjmB30RDBmKHNqQeXjI/VkQdKPt8Jv2pn7CaMCvo7Qo4ISijcZAIwdXiG
IaPTedBMG17k+PfIREcNqdCU1ntXe4w5y3GrfdL+etA8eeK0YV1T4MShteIoFeth1+Vvd4+MoDXj
kxp6ZeU+Mcg++iUjkfbD/CHe0VSa/KSgvhIuA+HpNEH8bb5TTgS+idM5W0Zv8ZKaD8Z9o+qkrPi1
Rao1jcy/Bk0MB503llQmhIy/DNUTnnmwuj6P9/LOlAwQZdJ9WUBPxUluw7X8tow0L3kIiHdymhmV
5e15Ii/MhdGh73fnU20zBGCDTuZZ5ULCZjaTOUG1PlzZ4cOfyYFjBm1dSdBQmovJmV9w4QPaCp29
wP4FIH9MvJ+BJzkEAcWiHqnBPxgi+hItcNdR0Isge5oK0SF2RxqQqERt+YhyKaRX40WdLqra6OFy
bnmhrKIzxOQAEnyaWdT0OHg99V5rWxQJkfHivCxFqRPQgjo4VBsun3OoE1tDaymowFZHW9Loi+L9
rKBA5zIa5KyVcDTqj4yLBX/bKCj3aTBJUhSGEdSjQNLYv93VZpLHmY0HdCoGmd6yqF8KaQBwBi34
1S/OJYXMQ2cx1yJWQWPzftISaVTrIt07k/Fj/SiVLaHD1sgURQ8KTojRXOt+7HwCuoeD2KKJq9c7
MZ+VL7InHDyUwN0AYurRbEpoKzGcf07zjm2nmPnmMqpDwa6bO1lBX+vTeH4gOA5EBbkZ3+UjB3yo
1yJnL7QmbP8FKAUif7K6oLP9yI4KEqjIj80S1JPGbvU0LS+HZ1tLicfrFSnziLfJyTfzQC2/ne2R
FTulrn+p8CEdEiY2UK4Yny+ycM7CvxsgH7sA0KzuxPsLKJ9uIPVpAjvVxAAjv3Nh6zVDPXcSUHXB
o0rSWrIRCWqodGxboMqykIWr6eDii9hCwxhdkVgrWE2/Nl55MRB0QiARthkny+bXjsfijJ1tgi2j
iXrJpeZvrAoF5TB81RMWHHz1T36SWxKVI62b8diekhv9QB1ka4Z3BFmqOAvK1UKA/ndaEsXYVIJt
fbSfhpw2KuYl7AuWBP4QOjtZRbp5efSQwparUu8PRuxXqKB0aT7DHClPalYCPbNcuFBJdy/IHs38
Ss/zh4DEENMFSl3uxkC+2m0t6tQp1r0giF+FhD2fhqQCFwmIDW8IHeUu7CS3okhZiSRWS4R/+074
IvWEay3+iAK7lUANY3EBqD0rlWaUy40nx3I+4BUtqvebdjeBBYkQeL5/9P1W47FLmtqKw1b40iQ9
3w1yJnQiwGQJMDpLGe76S9zQaOgX+a5pZ6KmqjGw+5PNsuHmQRDDi7BQRFtFwhiAFsKdZ9Ovs9k9
faTQjmmk7qmv4PJ7gPfcn/u5qNOfUiWtddEd1cFuhcOzCq0V5aw0ru4LuqIgLveM+t4Z6t+GjgtU
nesNGVrAlv9bSgeCxUoiO9tD+ZtpVZnwjDQPSz5nckt/G9AyIk39O+6secd83LMj7uLCCD9QdQNL
6T+bKoZb+O25hvBalhSViEsTr1XPUWD3yhz1bFoBcTMjO8IvYXJHeYtsbr8AmeQV5aS1luafaVzB
lIWMgxNh8F/Kz5cSuU87p+PI7h0cOtTAADO+9DCA3bF1JSr4AhIHb0sWOGh0kXEeVS5GU78K3dJV
NAaTuotFdLybqpV5a8RQvDXGYtHoXbuAWATbCg37cytmJhVi//rmtFneobS7AkMtlNR1HTzAJmDP
fE7r1wF75FHfmMXpQGuK06TBh58DxslNlk9MiJtcUJWSGzTkHBJDxsf+EKpdpCCCBE8eNDA0DKGr
oyYClEIBq1V1HAUaNZ+KgDSw5mR9EvZggizS2BZjU9pRTN3U6T9kFxDNstqJHkLsPaie8qugcut6
eyYb6EmL8FhVAFRK8/s0mEN9HhPj6GPHwxtasgTO/bBWOxUtiUfDAZ2dKMpzM150PPf9MIlcrLaR
5tXHrJbt3fqjimqGETOlIdSdZRc1QkMmCJnGD5ChU7UWc8TA1w0ZcyTfvBNfs9DVrDfjVpfRHUto
2z+iNwsixBAhJSszK7/5JcQvSiDmhoLhTB0NPQ/xv0Z8/7eaZskBEHVzwyBQmyLhViUoj59akLT4
/ZqP7acvveQ1lDogWAkBoFGaNpt2L2ONF8TRVsDdnmcMJqlnlx2kUm6zLA+fQEgWUB5jYUHkryfv
2gZ/mZKh23jyakdp8rNkUT/GdRIXAlMqpi++19hyS48QAZYS1BDtT1bKN1lcjCi4LADn48ND2mmF
iCtPRdqlmLIr+uJulJ0KYyjgQLQj2N9dVVZ7pOopoy87OA/R1M5R7wey2lynnqx5KYuRvu+0rceY
fNvyWKTkfFONOqwqtAGs15l2nS9MVsG8tLQh7fYpiRU7H+w4Bu4sT84EaGZ25GjOzmXZnVwRSpc+
+r9QBHmMbWXNuybuv+s7AGdzlfOLPITukYjb9wquEzkm4xUPoc0144Mbp+RYvmXRrkWaQKB91k8D
ddhFU1VOK5LnZMUh443/mo4CFVaGYMJ3aGZCF+J3r1FHwa0CSesh/La0Vth4s1bRdEZ4V3vMeMc9
3IhkJjuI3LT2DFG0qwHl/XX0FEK9Lwxvn/nNfJy0mMo6zK117SZbTOMqcw61NGPWTolj3OFUalXs
BMvN1UR1/sTwlVNJGqF+QayLBlZBBCpNCkJGqlmWBXMrTpBEt6QzCYGDTq3LeA+S7pyc29+zXhzM
0OnJi7Nhy/Ysy7SeaCyMqNTXsQIB3Cue+OGvZ8072JiN+KCkLG1/vLplIfN5vi1Y0qZ4FWsiA6f5
4+IjR0B1rfg+B8N/vj+rA4pRN9ogh8CXolCckYPiXUgQm50/ubLHApOB560vqd4m4XXlFk6FYc8h
6yP83TE0sNjWWM9T03EXBL4w/SLrT8LPEJcpiOfVLqj22k9SD7SA/LvtKam1lgW70pbKYWPhhenX
nb1vwO2HUhyYwcRlQL+YtHU6NH/B7qycXWLxlTNIrFi6mA4R7Qo8zOPdbV1tjGpnkWOvxmNlCDca
uRiH+LZlVVII4fps3DtggOVfJsTE/od6dsSn8Rf03s1cpEsw4ZuPO9Rm024SKTY1apE1kHU5wMCB
yV+zeG8UE7Vwd40Rv4QVhGY5u3bSofFF1YKWeSVVosGhG5DVy3LXTdx3Bj2NXB6AcfAfrGUC3wgj
IRAxhIoI6vlHET9KaCr5jm9VwM6z12LlHi1r8TkzHAa2XVR7w5be5Cp1IOK7/w/PXyv6+wnQZAcN
bZZO3mTXgb6vbn5yXHmXQr/Lk+feAjnNlOc+1BrgDktwN70bc5UKOs7cpwo85vpmlphQXWi4NvGV
ehW72NpTe+pxoGYoVAj1Jp+sxBev/YdJ8ORtkU1bCoT0oJtwalg+AYrzFVko3jsQuilVKDrwtrop
AbHIVdmOvZyFPYWp7hJarN1Ft+6glb4FJcJOdDTNZ46bwTqIU0LDg7zEWrxVEbtyr+3C6unNyou5
AVVv5X1NsQQlhfWs94cPtakG8mKOZ3hnrsz85ddhG1kG2UsuS0zjIFcnf+t2mkLEWfFJZ9Thrfuv
p+ghVLmGdtAOdnxSSphsNZ6lJPFqUxPYAEs0XxVoL/gu/XB0tsmDN7tCmUCsqnQ4siwZbiqVS5B0
ow3EXD5sZWXQjCSdoi1QEge21U0DClI2Fng4zWWzknjuGBeU5e2YF4YcxCmUqV5SPQsmihM71G8Z
6BYIS52CZeCkfJJWgolVpBcalVaXWO6YNd/0VJXrn8HG3lG+Qm247QSUCZAjhL1JMRx9w7SZSQe1
XN2qVguWZwOs1KoHV5QrXhZRejqQ6D0KIGjQDQyd1X36vqQfhDIo77aIAl6So4ZNmKPpcaQSzZ0+
axyy156MOgV4Q3jHQdUXOhVVVo4+1ZXRA3VOuxMlrmJBnaGquxbFNZduSB4lJcI+GezHA4FEf/8I
ZuNDtY34qQgsMO8ru4c+DqvH0bNEBzI68munjlKfH1uOcOkZaVTNasFusNLbRLJhJbjDzbNq5zLw
FIiy8Wdbj5flezOBJDegz9uk+SP+tGCyrZd8jnyo5VfOcNazxlQXlxh4IRhxz0J/KzYNWc2D0y9Z
4Mqd30zDSm8/tnkJxtmtm9ykpBlFc4dNbrHKzXK6Ibzoz36KE7nUbnR4bCtDr0W7SJptsOfLKFLq
XmvRrXFY2FPplx06rv4cTciTaZggIHlr2dGpBDUSc6QAG1kZ0PNw0uLjeo1nGSfH0M0NKJpSDl7W
OwdTLKd2i+37ffXN7vdjVSPdoIC2zKACrHNXQpF3XLsXH95Uy92MUQ15hA8jqCY7E81IqyHjrRvW
LfWhfv2PJfP7unNMkYjj+HcaEd/huu9DdkswzToL16+hr+TodySupHxQCJ8PotSeFKlr3XxwuVWq
EOEALWLEe+9CnArkbmLm6gF7b7/J8uZ5Msh8BDaoCNtUr1wMO07Mn+VFgvIoEzPuwpMET13+Ymr5
Km8JK0aX7eZWx80UVddU5b6KAvRngHqZV6sULZpxKpePNAN3BxicDf8LYkvdV+WIHtg3gLBJjPO2
CWJD0eHtMyDqbwQ6DZowSAeUNrtj8RiH/e9b/X5vd0/JuwKOMxWwCUOg+feXDVGcc2rOFscO7RFs
MDkkVtPRFCTydna9WS+5hRNFOwez+yRjyuW0x3d4MVY2qhvPgfOhgOd5SD8dyt8RGw9Hzs9RJ8M5
IWZR8uhMw/EthM14UjRGquGwKWQ74qcDCW463d8xVV4spydfzLOHF+RI4Sn/SICjbfgXGrq4B8fD
Q/amCpmzNPNPDvlncQHaZLMrTyV8htv36qIQQ5Hj269SmtJmxPV/4E54LP1XydlRGGrxEF75b+7T
ZjlweBci6Ge5dsOqlJDIeBemN/oFvSDyg/bZXwpRfz3gPoMCLKSEk6NGcoaUfSoaqZ2T/Xzc5t2/
sIFYhrLLMzCrkqdy+oUNr2h2fYbLErqRL0qfRiEm2nUf79emORujFbGfXCVmWTy/TsUcvbqPbD49
soD/tVJog2M4QPvzjft+nqLfUai4B+WTWCds564R20NvDVfP/n71nEAG6Id1FoCldOI4obHd8AOH
tN0SpCy69My4IjweDbL/4y2xEELIZ5RasXlqeKby0n9UXrDuPCDrHYDZsqckS464f1VXzquWsHqw
cy8aN4tzQFNiJEHI19FEcIvmfGHgKuQqRuQ0It/Qb1Mjtu0s+gqvqvGSTYeCQMhiRr2SfjomQ3h+
LFbYoLFMWV238Mtc7NxOFjJGiKGCdHxmUPn6wyQ5x7yLCRVunTQvPE7zzYmBcE+6kXHhtQECNHVB
JYHIaSKu65AQUtlNbCmMdiIMSVeb9SWT2PaVY/OqNBme5ZTfZZQ4smCPuwGzbYGk0a/nHC1LnxNV
N3gqrj/1EG6VRtEe396LVN5URJNNMqGSRxg/KPOfhWjBVezViC3vRDQaFIdauVLgWtuhT6Peqgtd
rjSfYaYDMJNTT5aCY0QhOScVRreSjjjKpwKTjhWpkJv2nA3fJ93pA/uD9JBvSJqnq21zlRZJKOKV
/5Trqyx74TIfknCHYyr1hmtb8LO3fViSQLTMcbs2x3M5KJzKW6ocgbT3p19+YegqxGL2ZTYi0W4s
ErMzfTn+AG9i8jN1g/oWkQ77B8EkwQaX62DTwzHktMtdduuDLUM8hFQblSklVmL+8sb1Qnx0IZ30
Ynh6hB2kuHLI88i3YnmyMdXUPpqM/KETR+3aN6iBgyc6kxaqmOi1Hk9dpoj+d1GT/HRkH6d/tVTe
QwxL81PMj8ynWC7CabRsWUgSQ0ab67DqFgVySH9jAlFMouBNki085CSuXnp4eNTG0m3khJZ0JmGV
xb1PElWtFz9T+UUC0Y5DekCD3gi9P54m+XnwLu7i2fjJvEdWKJmLZKWZwN0jzOwmWoMhaN7pjygQ
5reeuEOWrvHvuptB3Og/QIceyGZWYtwM7ROX+IozMb12pBcGPph/yyT7b0d+o2ZFFpIV0gy9SVpQ
Bxe6kMd/nhyTtkK6KNMO9ho4SvaN19mD0zXXjF9e9n8M9sgkoG3mUcdZAZ/jXS+C4O3xj80zKKM5
ZHaJiim0dVeWAtQG6oITUzs6MXY6O4ERT9Ngdc4DYyAN4758r6iFQ092EjAqEjSkqOMc9x1xGgBf
+1vTQhmZyV7m6r3yOI+slCksc5LkdU5+uxXaBG6R89S73GV9G0D1n+nwxnl5IzUZJO2mPcT+RN+n
iqYfb+g32lnP/rsO/048aOHi6J0egbvukcZPWNjB6BWBFiZYffhmQv38+9IVd6X0TMG7t4L+38Vk
qPmcvsoQ3YgS8tS8+kGgUmDNui0+2LnQxzgUYrJjHJlUx8vHXN1wt947UHtk5jp5g5XeNjp90bCT
VC50wKuKFSCXJUW6+BJjInVZiV2C1X09K5u3ZwFsh1azyf2HWn1twxODyPgfRhvAAtMlTUrxOa09
E3a6ILd2rz/AHV742xOb1YnzQQYzcEluH73gNN2BP3LGBlF46sSYki3eAM8E4qceWFpjzrfZtEtZ
9cYm2qc2I5em5S+dHRPjxepAH5kSijg/HSYBgPAJuGu61CEmsj4Eb21IKvzRd61opxGfBbVPdWSK
/cbpzocYkVZaTwdO9vtfsvvnMlYxGMr8hoMwW+alNFgoJiNpxDZyNln6CT7Q7vLpbZkEmyqX5bme
EK6PLO2M89YTBwOQFEPJDT84n0THf6wRx6b1cTRH6RgxqBAoMuM5cev1NL2Xkzh9ws3bYzb+XgtT
fFqa1jGfDUrcN/2UfLRCVrD9WFzaC915BlSNLc9rY0ws/HHStmcsOB4c8XNNezCt3CCqOwxTryDe
ybpaedjlL/qn3yn8XLFbrEP5pPTNAzFRS9bckuFOVgoqan6QxEEpIOni6llA9Vplh9u+cb6emIb3
Bidy07WDSxTVlE0QIo/M5DoDbEXkImAA1ocVz4nkB4xEabc40rxKSalnT+lfac2RKYgpjRQb9Mb7
9HChHy0Osc7+oIODx9cbs38VrvetKxIGln84hHATj/eJQFZeowbPbdEuToq5/4R29Lto6Tkg9tkh
VXhG/qV15T1tg+bOPT+MoBEZ9IxGddIYTPHm1kTyOGrV8oGkxIQV8BCxuJeXGpW8+VsO/Y7RabmJ
M4QuPbA90ZtVAxaBUTU694SW9X7k//d85u7aNwu3JUXXJRV86v4IfruBT7jVTm2ElOYUKXFOVTwD
AuDEKmN33bAI+aLf+tJBtT8d5simBXiiVgedP/h4RqVjn/uJKYtYvbXR1Mi1sBy1RMRBbJ718+WX
1V5VV78xZdo3pJupNF9bpqUS2A60F/olVy4tJrw45EiVaaDWg0UGeF4wGkzzrQlg9VrUG03B3y6w
Zk5U/YSFWzBpaiS1z6hdBXqbuPycQ7CTp/m7OSciJsoNehnz+86uueoewU9Oqfx55Y57/ti2ypoy
+QIk1Onha+zKYYo9FhOn+0rCKJtAKgQzKlvXsxMDkyRa6Rlh2nLOPKYU270KMuzTZ8hzM24gE44q
WHablSjkrKx5EOwgQ000IjZzzRrGl7nFCKIqUE91LMbxUAjgTe3pgSAGIakkOGAOppzL7jjOsIAT
/8/AZX/8YUOzk9ryTtOEHBQVQPstFmwe3yBrIzgyZ4JmrEieL/z/1tQLSfhpPAsrI5TjWGDXJ7Ks
KrIlhF8wKktBe3Dg5+HDX+LHlPqsIA3DZ0i7WRLG4xF7DueCT79YZF56a2al0O6XqBBC5Gwn23tY
9VNr5d1UJuqHZUqDHXoPlT9C9EcekF5hq9m34OX1Fw8f89zszM2gs+r6gX+GTeA9DHJGFuQ6AsNI
AZnG9Ao3O3p2smGGPov9UaqXbynrzVf3TjjgQxgDetAfxMXqPhkSG5O4kFuG5qNe/HNI7POfRaWg
8RXSgTaSjk5flYzLAJB/Cbf3/MiajKDsnHCELHwADMWqRVRuvdaC3bpYa3zn7hzwM/rEPivWSpJ+
so4UWLFli+sH7VeDUZeYhj+Mo8zTqbwJlVYYT2w5NEo6gOrf1yJ/mjz7pCryEYVj4MtVrqX8hVWY
FML58rJV0hpj24afZO/V2bCfslvXg6y2qywh5ydYCePGl6zWC7M0vsN6nsXnB4Xb7ndkfeNfcSJD
Nt8ec6iCZ7PkQpFqjvBBfexIsT1BRlM6Fz4w3o1/AgvdDpytvCHaxZFFaCDvibiK9l/A1PgTP5Yz
hu0ox6/c6ObcZOJpBk15IbnDUOhierNg0pOP77Zo17H8WKUcL9HBzuToNgpEczkjbpEckkmQBYCm
4ckrubpUCV2/zosDhCxJ2+qSZrmzMdyEbLjsfrUzXGNsIq3DomCNP1L8vIAT0ByRHbTXKIUcjEgw
NzEcdDl2Htc/RIOj7queR9OyCjIWEjUqGSXWMjOJD4GwZyHlToPJ6OM64VIkKg9gfUx9lIAplbmo
xrN5Dx0NKoCzBvKfCxeV0iFMah+Fwl/bnM+DA331FE2rQApFDhetL6e2aJIjjxDHNq1FfDV0h9W8
lkTYlQ3LaNFzdIaQNLNfAjZVWDChEGGfRXIiiL8fKwtCBr+GxqnZLtjzHlro1EwS7t64fXR+PLVv
lYP4ZUCJ6jGBHLdfL1aBCPfscrTSxlnpe7k7pJc0INzngXugo948AET7NLKtfLRWd7wgthndy8Rp
o+Xh4IuEBtE6Frx5LEJfbflbzMKAFkpWcp+62SxesZs4IuAN+ARA8Nam5N3oh54SRVxYePS480Iw
EDZ9KYTFuXD/mQtlMTygCxvQGQk96FJ+wDOy9klS6IFthMTR+63sSMLCqLnTG4ujTuQQKAMuQBbu
A7lHbuPlbNrRlId8JP1gQ9y31eePTH3Ipq32xM5rGCThB848jqJ07lfYWByUlfn641lxlZFESyow
aUeF4az4/jGrsS9fW9ndUBI+Dofug5VlsmKmVfYm5BAT1jkW8ypA9dBHnI6bj18Zx9JUZcmEDDGj
p8HH5I0zKKU+Myge29adkE4HM+0Dp9p05xiuP2haGQOEF3erDV87AMavLAe83L4Dc9gY7H0yOxMD
CAxtlstghawXXXLsVfHWlAORXsqJFDsdkaqACUm8Nwu8K99comG5120wHulNQj+CPhMBFHxyuSPT
qIyguUdZXMZ3DwY+9bFYcesP3Bsn83vysdEfc88YWDt/ZIq/67h09al1vl3hMEVq8qnxMxOQz/Lm
TQNwDFoQVzGDud/jCzia6HYUtT/fE7ldsa4fWFp5S4XVRtxSSm7xQG0GdtE4lvTOvf9aYvORjbtE
08Pp8LEVdfVRB/rj3+AMDP4eL+y9LN9TnLel2Vi5lsMnV3GZMmRdo35x9T0xyHOhol67p1mN1mm1
UmqP6T1cBIDZXj+HWQ2WkCV7c5xbxrU1SAFRfCkNHAz2uxVk6pgIiU9B1sdn8CvWfiHFpa36mzUM
iE5oaQvkcxJqkqV7g4cAaBsg29YNLNreqqlR9/ou0hpF6uTagKCToFR5Qj7lrbgJz6FX8s//THM/
q7Tj9AySm7Tga+5qDeHlMSfKJNp4UPRxGgrDdFlZ3qcH75GB/UmiCpMKUd/3fw8Mii7lUed/1Zpb
YVGS5H45OWVI2TVBwdeCd4ILKV09xAMKmS2jUmoOGjErThFWXsWAb4dPOKBISTUz2HdWyIwHdWVO
QWx9kMl3CiCDmI/t+0RS+iHO1ysXh57UI787bAm1gaswRkeQyjWh5KaPf3kHd0LP8zbBrZF+4AoG
85X5wYZr9eqvOf3iB9DiA82skqYzzApTEUhh4SGnHyr4qpuBidAlBCYDU0wTw/QFa8XmELmBLp9f
9GFVDGPpiCCrfw7adCPWGZZVhFZLTA5BsDRfnRskN4FSff/jKh98XyrkEpUwzq0Ofb0ty7rAZsm0
xrqOacknr1Ah4sARy6DmyQqDGSdmJTe/MAyyqukKB2pS162x3Vtq2AzLrm/lyuf95HaWcyHC3d3n
HzHB4tkze0ci4Gism6mefFOr9TjEWW2bbEJ8QjNBGNQdvAY66+rEa0rf2uyIrUysCoCAZ4ZCw/d3
jPDpxOGYyDIUBrEyT6g7Cc1P+nPPxH5NZXWNuAkqecc1sXHv78P8dyWAg6ithAaY0OGYNYWUnEza
oookLdadK0fbq80DWELo2p40ouU526RjaTF+zJkHmGYHoK3A1gEyC6ewFABnLoIOwnY/HKKtZMCp
aozEuDfu18l4mq+9JqUHwT+H5a8TfqMedzP+GdOPf8uBSDxZ3KvAlnrzTYGXhGgfzKY/+sKkKvyC
Vx+YDhmnrtyG34MrsUjKWriRbyTCQvJdji7W3aRwatLiuGlnaZv79VvLI7CYZP7cMbjH4w1aJiKe
sQhImZykhuUnabgpkAkmBjMfCg4AVeemACPhqGSr2G/lJOyi3l1Vay9E8YOGxOFma5g4xaEy7Lhk
C1ol000XGa1s0rtdeVW3UQ8kaELxFQmoHCXbBZqF32E8hiUTTGFXEMv/Z2pTdKAzrbbGjX0DO7NV
6oVYKdI0ISXY9HVH+NZRrLmfDSPzzB0E4m8tTquGSZ/qmNYhj2wQIK0XaRlCWKc0q0yXkV4lo7IG
ioDsrbk3mV56oh0jtUYdyzbEO1jdhGgMajk6bBjp8D7e/2oGqfnxCnipLFCSUkuPiFSfKRSluO3Y
CWDO4Yd3RrABbMMJaod6hs125Iy3zTF9+xeP89smYyf4LGolS4O2WA9NAGWRStb66EB06PGNJNvT
sFk6KSrs+LWnjs1+Y/Z/K0MkqfkTJFWf8TKTJBKaGv3YXYPVaAyp1vNRI2gn9Gq8h8oZxSWV7L9H
jOJ86FANc2G3hbjiApJk8Jwc5lLPfV+AF4WHxlXVlkkmpyHDnybBGABMUZoiwIPNWslNfCHWR+Hg
sdq0Ae4LiUNtc+onX0wYzIKzJ/kmM3W50l73u/DMa7b7njZggGqGrUXLfeN8mzb/AclrfARlvQWt
WxXMcPJ4pGHHPDxk/Afx1Rx38rElhldFN6YoHEJgmz+TU5RIG5f5GW/U1GOH9DX3VYX+mEa1B/OE
0ggqY0UXyJkPcCd+hClk4Qys2yM/MM7ChEiYD24HBXUCaNjKxlCKGmO2/AhAQZlmkvmSUk8677Zq
fxmIjlYZSvHhXc/PegOyuavwAnlpegXMOQdinYWhOVt+AYND5Zteo9ELYHi+5kIsZxl7mYztDz6t
VVXnQ8z5MF/ZLTMjJCe0p82Q0h1Q2nU919KIgKofO9s0KWR9TnDcst2spZK2P0NYkyL96Re2a6WH
kSTebmA0lYivfBeXMKDOKS3HgrEFOYnKW6kgMtJEEMUFRNXYtEbAwj5Cnb2y9Y9eeMbVcde+5KhP
kdOGhCozi9t3mMdUT61YiJ90Vnf0b03wMy8ZFMHKqsoTtyimbpjvEtanfrXGRBnCWyqQ+1yOJ172
voLzuRKGQTE3uIuLbE1gBo4xGX2o/3rwiKglY3P/2tuiJzUId0CAVhR9kiB/8CuVfXBHMJr2VlF6
0KTqVsMamBPmRW+INm+0+DnYdkNXE49BwQvLuIyyKyxUmbDX/iHAMgw9gel371Nyxzmi5vacLPDz
YFA8Ub72VrcXQLL96NIc4Kr7iwnKS79FJ6wCz7ugizPGJUhK3Am6Gbdz/N3ac6M0P+NNSe7zmYMI
+cN73XeeoiNH6WNxxsE9wnrUriYsx8GToQUw6dUBgKviisJL5Y31jUHKGGih2th0D74nyDjkV6sJ
JTR64YG7+6goRXFHv1Vmt2tknzDmgezopV+J5FXDrzxgexYXXbr40qIGfi+VbTpVWFNBvpCWXeOL
2qKUjKTeNZljpoNuVz6fQKRI9Rl+zM4ZutebZawwhBqHbxiG09+SqoqMU63QGHvtnRNZrvkyEgAR
UDzAG8AaRhieHNzogt62do+yDGi9G9/I003GaRX3kLMYdoBZu5eyK1vPyZeHm1WTvSLkcmPi9hA6
PAxMvdTxptl31pSDxoSlOfZkCGX8hWqg5swd8GAvOwBuzbtEUQ9yO0pZgVOKSwOcLr/t9TLr6zuE
ayLYEugr0Cr+mhbxY2WiG2lyhr9N6yq9L37IV2SyE/CSv+xitRJyVsEQnEBLIm/hMqDlvOcR7VQE
+DGIE/QF8YzPTxN1cP2UY/0PW5+haVpT8b1IJGbUDy6yZaNExQP/wffrlHpNZ5F/bjO9VwO4Z8cR
MmtEUtXzqFukPA2inynu+H91mwNdLLSb/NDRjIshBma/eH41I3iqSNuAZgtNzkJGKtlZLIUKc0qe
ksRXyZ+IyqENdsxXb2kE5Re4XhMRNRbGesv+oo1a9eGnYv0nmbB1957YK77etG2GLFWtIr8SbV0W
nsjUYBQWdGm+B71sW5Gy+bczC2I4ADfJMsajlneIqHl0SSSF7a21dL5VrDy87CvCpic1gKieJ2Aj
IJSXjHu8OpurVGr3mdCBCANsGLcypPAXbmnwaVXemBz0kN0ymY4aXLDWxgtiNcNBNpe1IqAxen8a
EHyEVqNLiknCJ1VbIcDnjjoiGX2BTr9sTcExwEcDa8htNPiv6NojzBWQvsaQ9RFveOpUWwIL8zBo
99JkzISkvW3EFLEaApmlm5GObnF36Ky1dkUqCUVz1rjUjmMvdcU/puO0H+dpfmFrIbIhBZJUKsly
UKE/sInClzVkMbUI5sr1aMbUGTP5iDRL47BtakgoGz6RQzoM37hbTKrNz4SZuaWma7C8uWig5IWd
EV2EQjVVVX6SszoNWLGWVoOGftcZoTf/INHA+ai1tkpI+AnIZCq6CE6N/4jEVVkr7Sx5oaZxX5+j
NdneCNW0w11iWB6E+SthrgPbAyOqXs0ajT4FNhKV4NGi31L8tu0IhwHN9VpM0CUuvAp8ci/fvHQ9
PMz3WpgeXjoWdGcGTMqDnp2BZctx7k9f4RzGmJF/Mx6aiuNXtfKztcM/oXzBaflq2fBZgSJhCprP
lpjuUAqZFghqCk5d3BZmE6QUSenh93jj6ESUTJ2ZRt6t3t4MZvGfcEhiZPn0AV7/WxjYa++tMmjm
Swm9g/Z5ODf2Fc0IlktOVMoahC4ajltk47DvCpjlnf/YHOXd+pGeehpe/3FJEZH0NgMsL9YS4it0
WzeAgH+5NpSNLzLDNHNniSf2VAiyMSWOfC/WcNeMPjnyBa3xwW3lkPfgfGR/kta8DYdV85BGzAf5
Hrts9Dnqd6k9hPP1VVi5pRYtRaJeE3GlkGTKNVSviUJ2mNqNn9ayImplxBTwsD0mro5BK/kA2CKR
fKWFJUWtCqiISZZKSWuIi1+VFsklLZOSSV1jYKALMrmgPnDNHWbnWsScp7a3xV7VhQTY/Y31p3dJ
KWhxlx4jyaLSqvKMTCpUxDwsoFBXjA5C7uH7SlrOj+GsPuaQWf6nmffJ/ABLtwvJGFBeDKEb8Bqp
nk7T+QjrIk2pWHp6AhwGSnyLe1Y+Rmjwk1GTaSErN6DBcSrwLmRCGTrvqL1G875iGCQLx+RI0hW3
9BEqfYR0gzGYZnLri8Mrb4H9NtHKSSpUynq0nCGVaOzccRxlIXbFMCvCaRxWL1TV60pbSGAxDKva
UsTvdk2cUUn3khxFjd8rulMtv191/ry+Qt9oV0BrBGKmw0o0v6ZEoEfq5EwtoDFmCjwjnZuuQ7yv
IEKGGnhrPCQQ8BbuKhTuFP5UPeRukJeXlr6IvTdW9kyX4ISPGO+9NefELAfAHJ8D4EPzidxrWw6D
s3pxAxZaBaAY42fvQPbvhvtIz8nGfBmb08SILoEV2Xnq5HznoEZPkmy9dWFlUr7jmnLlkzOtb50x
0PalwbyY2KxNleKXNncB7uO7qn7Ff5oRd+VodvRZKzKNDqxjTOrtu6fuvy1eKHzPM/C4jFR8A3qD
EDo7G/Cvp1o4DqEGNvhx0+GxPDG7ARrXWLGQDpumpLCqQb/1sWV4zaHUEiFnuxTDCw3OhrJMyhoi
OWYUHcuFOyvp23xqxw/Tmbxdum/4fg/gLPN9qCdfRo65Jr0/ZlBh4cdw5o6xDyxEG3+psY6u+c10
/MFxbMipW5yKCAKEZFhT1mEyM0S4RKXxoHzdCvSFEzu4hAKPAwJGdichPZPHPAfwYSk3aXwswSmL
LZfmaa46eSjntBiboD/OKdQOmBq3vPWIhSJmlZDC7zZQPIWoQOJXjX8/dqJJGxmXjp2fyiqVJpLY
cuUN2S9brfxXj4GCSJKhniPUFRbvvOslhui+Qa69SWxdblx9AUKKmrPzSjYK9bsOu50h2QdSZ570
V+oJwXmUkqgjQaSYrS1d6FOXN8czNPhYPK/lDJIKvduoHI3kaozxq64AmrxOpMNiPdjfgSVstHbp
Qk2Jle62Q3I2C0kIYshxvCDBs1Le9tckPeOH09clD7F41R58G7bt5AkK7DvuFPf6L4Fk+x8MHhcz
ACA2f3K2LwNcUgkcQSOzxT9vZd6YvugN0yDTnihf6RjhLqpUpONtPPTuZlAMFIIR0pj7oHntyJHR
relDhcAMr5TQ0PhzuqeGjdYeSJPesACW/KjHqlbxlMZjAgJfozYgB5Ib+jtjp4EwFQuBNAFHCw0Q
Mpjv6F/1C5N2BOALfel/hcX/Pk7zug4bIBFfjInEYzZFJucW7XewAaE11YHPcCi1GYvJNOrBVFiP
Wiz1FLnSKLwIhGI3WnMjh+Xgsf0rPmwfAshA5p3SUPhf+7FHxhjf8mzanpIkp4s3+66BccZdbKlO
L4/wh7u17Jg8kDCfTqp0qrWdftcVDQApOjNqS3t53YOoohPJePME1P2++kBTQBYh4EFPONU//2fx
LdfV4NPRbMK/CDEF4gVOpO6aL3dRkRFz7Q95gtTmIzqFv0dUg++tWzcoyOyzIzaEF7lTlyk5SP/M
3OYl9fsQqnlucGywAtCsV54ZbJZCZagKQW6qO/BmgW+DCxJ/2RMxZSC/VayctLZIXZsgKySooOm3
PIph1ZxfG7tLjiTlEH9yZgevqka0RKQ15Nv5GyLrLdgaVXja7dtPcakNcu576b0UYF/sCtd6u3jZ
P6fX/+wytgKlaxJcIhVM8qoHGJ0Nj9NKP8MflKAs8GFhkxGsIiTCxYf+76/euIzBoK0C7UY8Y77O
7Brcg4EreDf8JcACzaARg2UUxale1O30VOQxB6g0enTeHlR2m+EekNp+BLl6LzGmOujizp2p3ttA
se2Oy8qlmU5W1zcp0Yg98kT3kckCrZZBdoWNUWbcPiUiK8lpNthp9Mt5uFCM70KrNFvpGH24OZ/M
eZuLGmPq+hdXNFPm1SSYHm76gnkk+sK/rL8VYzB6P777MztPytgczi4kxU5wCmSY7TubOAWXsbtF
LY8lpGc2nhXFGqBsF86J1MWp1joaNluCtmyn8lmuVTHIRPlAFIGug13J1hnVnPUYID7B4TdrLUhp
/IGLx3J+dN/It0Vv8uHhdF3bYJSvOs5B1cEDcrKwsK8a3G89zo6VK02VwbR4p8LDEkewnY7EFJ7n
uKx46p6Biyg6dgLu/db2wFaH7EvnEt6QmxI3dAhdxGKwN8VJlJnLq2A2N7XVYXAI0AHKnMVitvDW
b9KVWztFAN+uQbI3lHqSmeKS9kEQ5KQmqmmL7SkGgr8mD5RIYLG9ZKUSVE8wFfRPPJJS3m71QfG6
EuqW9vjclIbHiN6G6DmfUgLl7fylJA/bD98Q7sl8rAFnsxeRLiN6202hJ+UoFpnB1R7RI+fhij+D
u8IhKJKyRKJ4YVkaUBramHWe04SMZjJi4dtmp4PqGOGvHkJ81lvvduwJNk8CkDMra/QzXbB8HcTu
HpGSYfi5V9eOHG05iBRYhUIXycpEUaXOGWUtj3XdVs7UCIwnQjX1MghHxBQIYP0dFht5HEm/cLtK
3aXniZ29cJmd6sPHQ9rpPTCZ8P6udQ4bJR9mlTGXjTl2yFYDt6mpBdmaWOsWkIubkcUWhNs683Q6
HlbZA+YZdyLZ0fa7xYTj5Iduqtu4Qe4E4VQsv0LrbqFwYfMxZjGw+QOu9By5MKlNoUEePXOnSSP4
+ih1Bj0TisWmQlXcO9ckQNs8FZLSTapFCDQn+N2VlT5yi5GW/tEn2To5AYf2GVf3syMj0CUsKQXd
+1KOnJHkYfImhZye8HMyGfzF6mIWmdzPSVfnhQyFqPN06ytpmzbxgEEGc2nhTcCTqqIANOCGbHky
3a69dcx81ke2xtzYv3SJ5GMLVOkcsRkpXfCddbhtP4KS4Hv/p+TV2GcnqKmzUrCdZmkHwFhRr2cf
6mvX/zaRBclMtnXlGis5v3TdkmTt1WZuyw1YHL5JWjwLC9ai+0PVtwB447Vdbhn9FKRCyDm/CmK4
Napz0LTp8ewYw01yJCuMC4ZWfiT++zHRPv+/YGpSwKFyNXRpPf5poWkaFg8Dr2G9Q4+haS2xrtkF
oDmyH1iol2tqMMKZObqVr+8XSeMpUr8HDcIG/41eS4X0fFccS3Ce39F9koyWz1kzgQRlnTbycKLk
7RSsshepKKYPS8SZ2FE/A+kkuA+VtY1NC6uRenJ+cx3Ox4zdlRO4BLPbHr2RfCRLEV1MI/4KHD/f
dSxVokXbPH93BKV73+ORg5f3lrGHNbJWqaqGX9l54Ak5e3tJCrEGCETmmaJny+mC6UI9YM7kenEu
NaJvUflVfKH3IQG8x57kVJoKDPFzQsC8CzYflF+D+qJOjGb+9G0TVQwTlI1QKQ+E74HelCX4cj5X
v/nCLwGyNE4mdh7AcvJExyrep2PoqmOMTBc2dBD8u7DSUdkK7ohIV/E9uJjIDanzPTAu54dADXTa
K8ZNiP/UZXvfYv6KRruShCn+KHg11QaNxJa9GW+6UxjYNlAT2pnjVDh0p8bFv6+xUbko4Z9gQQnv
t0piiAWkAs3WotKE5v+JnAedOUacmorJp7RKK1wGGioQcSNq6UTxsmncvUdWmn+/HNgbeKTT4auY
WcxTaxettZ15BWn8VPlbdGlE+PkShZXq9xWFmBrrw/L9oLbqIbBNv9Oie8XawkPOC2aPv/DkosbW
PnNDPWZkZp5ly1hoKw0/zm4p9ICMnXurXY2CsZ9SCmIoRklhNUv4nONNVrfnwuVaajVNM7WwqqkT
tzb37k14ePJTkbCaVhK+T1Y1MbAQMH0gSeWeRAbYjvcThlhnpBi9k4+P51y9u4xQuO1EO2k8CcI2
V4VIb5qslN2dMFVlx4/how/135pHSnmBj2i8XSxuwHjMsuQp6giBmvNbvwWinunkSbgzDWguQjtR
DiPpzgKEOM4kLD7J99P81CR+sqez9cd3bC1ayaEYLobdHeib0qu6mG3CRZj6+jDZZkvHIPcDC3Zs
kzbA8PRhBTNl8mrTRIdOzMFIokO7N2yRNA/JWs8NvSkwuJU5dDuE/Jfvb7SlqPwZ66Yxd5IPPbpm
doUu7W9yuM6nve1e18HMCYT/m1czsbs9KGzKptHq9Si2vHdUefK2Rv1YLilDQuUL7EhV74R0EhCW
gPIUzm6EC24FUluEyK6h8K+sXvn5NzdZRV54KXAHEZ8bU5ejq6AwFFeZRdK1ezf0WSSXno4i7t4v
zbloJ7jJ7os7LhUJmBCW18uSLrAX7LkyX1sPqyEjgEK6n/gqnmlgnEsgIOha4kTiK4cOualub7Lo
EprvmbQxKfbRf7NL1+lrNjGH0x+exf/beC73AVhWAARtaSayMQfJCm79sn/nHK/HHlXe0rlGTBWv
gkgpr/tz0i0fnGsDY5dnAuZlLmbbEtHX9ymb/TZMbL4kxAVMiSUeUa5ZiIcrHsMERkCTHEYy6oMF
DtHdZV4rHMDPtiHXl9myjSCL1cnUt0SWbTyYjz9YEaZuvVcDcrGxAGwt2Z6jEIEcgYIlhNUJxCOF
PE5HU/U1KpxKKTwBHW04SWYdHrlP4EDMMYBxOmgk4ArZa4OhROuHxvP8vlX5+vhYWfqPsyk+whec
DpfAvTXqthjwc7ShKHzYoT6v0Qj/2boRu8e1d7sfX94QjN9CI02lTu5iC32VE+LqhXg9yrO/lxj9
IbdIpiXC+sxqgfn99a2vlzuldZzQQY1knzEyG0etVXQ1cd6Fp9Fz1LdFQ4ph5C/qPS8kb3islEwa
52m9+IcgtA3NVb6gAABpWQdW/13S0rCRrfrTm5ZJCQsiL5sE6zX7KTIbKBPRFx/hrjS4ImUVULxI
IZEFb6agVDYZzOAoce+hE+TbswP1XZTqxCZnoKvv4TqtI/9y1jGvIbDVDEcM3w6QpVRW9bCPuMRs
G8t9oEDB0T53WqROdin5nOpg04SJJLN5CZ8OQW9N8/UWZyP3WBH/uA6ZKVA0vz6vr+sdmQchjuDF
UsM4WsY/TBjXokC00WZfssQ6TTgUEKGGCLzla1f//Jv6bv7rc8FFqNmptlfw73y7WvgDiieZRqgt
lN8nxp/G0eZJjg2r4mqIXMkAPgdEq/x2MmBv0LoRo4oOnuUzrXJ5n1TRGOKZEYIt97Bz1whWvnwU
xOUyv5AEt0CroEJYXdKk/OcdPkYPlwfD1pRTK4P9pwRTr9CeKZ2yyGH7oPCVBphDAYxUW2ptbrs1
YvClNTKy5DE1HNWA2Eil0znclI/npQDmeGGi+UhNT8z2pcMVRU5H5sHheoSwBV2CRCZdRXt4KdBu
1u0HuwuP3gH/MydPK3dzfS9KTL4KgEf7CNhMhKh5pF+uOhh2uyixnQwyCY7K2mc5uYRc3XHHMFvv
i5MJZFLNhxqDDTy3Oscxy5UDWxTidsPC/hpI25HlNKXqs0i5qhhQ5tMB1HrkmfHT6F7tUX7mG7az
zDs//dsiV67F7bWe9HoyOrOP6D2z2TSRtzVtsFzRX344uU0PCEXX8cKzuw21w5rlzO6EEJbmfiZ7
f/NzrKD2+mVLVJR/cndVEIFq5OIn5RElL2nwMFQ39DHUaAQ1pL1XnGXzQmC9I9KNCtD/hyHytkiy
qn3O89CvEZd/sqE6qWK2pmb3eK87Uo7El2ircwweh/ZxEXbP1LstDsjC6qJwQbR9u5UZtFCDzgpd
gSAHJFdf+9buUyHaRjyVD9FsJ2aUHnlYPT22zJRIZOvxysZyBfQwy+F0qxlfeXSERlcEna4v3aZU
Egb5mkwvgYukRpW3g5+/2yLpzA50MsDEW+nY6wtPzSQ+ZCk/Ph3YYRqkgvkWwY4N6CHa2fYeVkDl
1orcJXrd0igmxuwIUcN7DH86BLyBaR8XeJ6L44y/ymGQj1CmHfxQS1na3P+ko4kP8g0OSCkWiqg/
OebLSoeFNvegcS3swLTHj+zr243KCyjtw7dqC46HEi4fHxRJJlGOh82jhbR2tewPMJ6LWemU950I
p7mN+X39FCym9POUqvpnlP0g6uxPv2jbbd/wokJKnUX1RYGDmf7AwBML5KEchArr5NAY1JFREjXT
QDrfSev6cfH5kB+lHpb9OZv5TRy9zrxl89+JWjKMfU9p/zD7rrSqIBPM6SZzwLorqVfRwwQPBge2
A+j/E/CKY5h/Am9jg64RVGyirnfCLLHrEipinO/5zRwKNU4CSilW3QvQL//aWYzttPV5aRavP07B
nl0uMtGNT5vYP8Cat8JZkZy31DEE19VP3tc+FjiJLFTeX9JU3RobGyXUUGNrgt3syr5VtdDdQpyk
t3SKEHMxF5s6uMd7vo+nj6DGjErOPHYnexMyT2rymUh+a7pJxPPISe6i9m8gbUcal28+tAc0QbaJ
dokkgJ8SgZWOf2GRPUcIRnB6BPiG4CwFdEQ85u9Dcgnlirag7t+xKKshIz0kmBhLljhEvU6AszHT
cNuqA5bUp7xxC3/Gk6qwC+eXyLbIFJ+MHoB2JfxG+3EQQjuwVWq2pdDVUJmWnTnKWWVYGvspdIG2
ZkbJldNwjU84VH6+TeawnOTG+cwePUJbhCsYMkRJz9SsHl8wS1MXZtCXwZNLDyDDyubOrtK3qsMg
la3t1CGXlOScls3xCp/Hg05VS/Vw2bPGN+gqvShGaddJd18paTUwEztWJCqBqWvlleZTdHAZ66eP
V9r7w4HOC2Oh/gM8GVL1ND8szgdESaWil2wuyOXKsDOgABjQPQTdHVUQbBzaawbZPb+aUjfPaxHq
daUvMyuCVkvLnrsVMVgUNz+VXbbq1sUGji824q2+p/BJjoMEZoLahTq70d1vPG68OQsTO097UXcD
lwC54/OLtotb7c6GO7PAH+uGvQ0Bxh84loNsegOmg+jZ717x7auJi2V5RVofXv8fPEYnUm6c/F+Y
F85LcWc0nNpf2brsBkY7yD2SG0MBkSUjty+38gxra1aSAyQZ62xW71+T5JPYsTQ73p2PjIi6kwMd
kKCTXnZff+XfGprBiwoYhJTclE9JeEQcZQAn1mS73Bsyv5VAWqIi0NRSJH1kclpkC6BJLR9t3qmU
gH3Z8S9VkzemXIP7P6MvCrN1g8BHIXYQzDsPkYxemymYvitZqbJIXeRQiYjWPD7l47ztyFuJ0NTN
vD3ghbdhZEvkBR2kZEr0aOBXVUrffzDz7IXHCSu67Em/BdHpVTTSsrP44WxnsB2XI9k5aP7fOTrR
hw1w9jmFqj8LLSVd+vzTtP338K8SNN589ceJ/BqWYxHFbtujbuhB7AUy2g7yOQ4DcYvyYV7YOvWR
CcNgzkYBlVxIpArRNDpDFb2EirAlK5LyulWEy+DBIFRbVUeAADFJzx+nnPBpJkPsHM4cddg8Q/NG
frDeoxlEZ6F/OIbcziHv0TEbYwdKjfsk4Ej78/VMzHN/V3XxRPzhTBGmdyds1MAKjPoHi8+eHzEv
VH6FiS+dJGzWBX4JC5fdkK6msx4vqYX0g5OzsDlZ2gs0BlbCQcpKt8a6XzWtG9JfjWqfkSl2swE/
QK847OsgdGhC//eW871Viem4M2BVz8oFHFmnk7od6QW2BPCQTt4qdLDrieT5MnK1k1CzP1cc0Bba
AzK/fcSpEpscZhiyUVORGDxqx81lZsF05nw0o5GSYFXy1gB/CYF2/0uTRk8apIFoRZRLine6qUic
05hDS//ffMR7ZcCzIhys3fQ4FNQVLL1gO0CdqV63WMZnTkbSKv6WJ0/TTZijuS5Za0joocoywd7o
EhXUclWWeoNMKmowhShpdB97CLPjWclqmK4k4NoOIGAjHX5X+NaePAkE0pr/XKuddgOmRyJSpww2
WCpwSI2z9KvBkfFZmXhdyWri2YAZqGKfjee7xQVrDvEIfv2+rNj4kEbrb4YxkVXP+pqtYsU7pMwr
eqLD0vYPZ+OjYrylVuLcgJQugasNwbLT+8x9ElccbQkqLdam+rGY2ii4QXKj9efzdevLFun3+X9D
bk9lDn9VIZxdwWtuteroirDEu/J5t/QwvhRVK7F6P3wOv1SSsYiE32meSykaCapJD5QKWnxK9l/4
IgtIFAPznx+L/nMImiPPzgbufsWFnwvJMqZBD+Swd3/t60qq8g+CGB6XWNnr7H+Ihjz8yRT+jDKV
7JAeqesq2W4o+AJ37tt61IOtf1j+/Y01xNXi9QGWSmuYGEDR/8feh66LxlIcfpxFSpKUSieWwgZr
9omD/LfpAQUSWRaLk2ZRLSO+AiEWAk62HKrWAdThblDOM7O32WR3jiT03ftJtPPsMyZsPe7fGlez
+6Q4w+gTeqjFpB4Gga9kGcnpvIDa8M+P0z0jEduAXaPx59BO10unq0+05o2XPv2RTlqgK1mW/krm
ImDRWziAsU99oTM4iJcZQFnK1KQMHSqM3/JuA251EB7n6P/97Kc88juZIwivASHxZTqnPH+iXHL1
Bmh/i0x5q4edjnsLz7RTQ0WkH9cTnvFlXLor2b8uyuWpMmBocaHD2+ucUmgqF4T5CYO8DkUW47uW
npYEcF1mE8BbcAdtI5gVhMpet9OrLAz6N1hpwzHtwuO0hOH3ets3FW1fsBKrzCKfCQBi0oOdVH2E
GK0M0pefYxz78sgmFtuGQyatASB+c3XIo4Iy/XJHuJlVi25ywqV/mqxhn2Z4TpXRGY8uiDcxcLne
n4yVX6sEk4PItWeyyEJzrLoWJb5xXWYIMagxqK3SjdYX3LgcSHbmtDAV2/e4+uK+0ljaTK7pqiFu
RSNE4CSz7dgsc0zD3YA4JRmLdw2wcWWVD3EWlo5te2zuaDWgQZlPqaQjWh6Oj6pNRXbq9VUhYNUm
5s7Of/5dsSaxtFDBHl0CLS/fsguK5pLMDNSw7IMNvH7UDrhCuqVlK93QRQKfcXTeTswQwEGKghbg
W1eaGmGioEK7LK4LnHs8PPKKDMIrSDE5CJhrmV2QAIbOoQpnrXjjhubQmLLuJn0aTsb3/xHW7dEN
qC1jI+5q2++ZemfpWVYvj+XJvo7qK5De+/wUYmQIKjde5BVbA12dG1kYrECjDANVCYIBsOXcO9+j
5sMqXbrdyOAmi5dsQm5L7eQt4yggt3Sew2j+Ih5VcPZWleNCbdS5nPqKnXXpsfOCA+hSNDlMVxK+
8wuXf0Ir0/CB0Jzj/Qoy2VYEgpx4Us9mYvwdwORosJX/AChDVpJgxf1UxkOF7WR8qTZzHAo12NKA
ibweP1g+e9Ge4DRPYW6Cw2U6EJDrejWAsrc6wNMUhpjqa5bq5whsQ2cFAzHvAyQ1U129dQklfjNT
tsayNpHgsDBd5SjeNMRPPwzJdze0KP87riNRa3DMnAIv8SnQ2SAwxwWwyvjWtaiUMwc070TUB+29
Hr0UmFrUHkiWnu90OdOkYF2HfRyijemIv2Q3vE3ajwHaIZsqLM7Ryj0mMsDOtGEU11xZJcjkdeCw
59weg1MJPKjUpLA8Ia5Gwq+1espBXG3owbxXGOxBrdOIyAHe9Wnx8i1wef+cLU8GXXCtZr/OgDsp
/s7//qujNiv2VC90G+pvGe7EAbRgd3fvc3Gzigpo8E/SdYSKMK3GeQbfEk3/aSVoFlaetR6b2qoK
lH5T4b7TVF3G9u9jye7J/Ghi3FhNNP7L8QdKawQqbtwdBcS7Hrnf5Mtk2DiSZY4bh21DvCIBEq1g
heVIU/n5rbSluLJvL2C6mvBxb4h8dTGT+YzHfQo80rcAJZiRJ8eDJ2bj2bsKYsvXTRHmGyO9+TXt
iEWmNfDpCVA1KmOxrbpH9UtO5g4QJjOZxczKPGnDqQ1ievFD40J0sRiBqzVGKqCMl4LPV8ckwINs
FEGWYH+IC3mzZahm2VxvXjoadpEFIXuVNmKqA/6qT07tnJjX4EIHgrnz6YZ4h0x1YcDmO9rDflJs
ZSfQgH4eUkaJ8PN6AZSp9jrFrvBgZvqbedGSYZ8khwh18U0uY2D7WxZ18aE0Y24qMz6C6FjUIKlv
L2kWUp2nAjUky0lZEV2wdKxxU8KTdsTwe2SVHLzoV5ctk4Hy8GmchGNd2P/dmiyEk7a/2m3LgSzl
xWmxiLk8ucfPaFjhQ0oK311FBW+T7g6ZvMQ9FfDVszUIMS6KCyUjaBZFRV5uzQsnHyljhjaFWoUC
RlSBp+tL2mhFKYAwpqt9baZjgzOF2YhNKUX3IFcIcecpIApKQAoK+duswONMSVHLoIqKRCE9pjUA
sKPnlQeG35Ob/Ra40j8CSj85FUODUrIVjxY9niMxeAtIVMYq2Ol7UuBZSXT/44MIogTKdVUEKd0D
EjIxPKiYL+UU05mVKOY0YtfSC/8gPf6pNRyXSvi992JNKYJ7ozi01UoWp84EciBzeKwLFvNPMYrj
TiwXKVMhP1z783N1nSZUbBzFVxTnPwmj4IADXicFxxhrnD8ltagaANpPHwyRxAA+lR7Y4uYxPzv2
80WD1IwWjGoO6fqUHTvsGiJZvtEXuZbN5yFaGvF2vQWgHS4YhTN0LOmLsCFkmf0wTwDX6jGoK0yw
1JwltGj2GUxtdInwSSR91MCl6XWrWMZ9IiTMuIiPPEtYvIV+9MZSPbbl1RdyOtyb52Z4EG+f6Ocp
QTC/N1rkxkFScPS1UxEsGxNv5hVqH5Pj061TI/rRMrx2poJDbx6SUeWQ4PqGBEY1CFxsr2g+oDIT
f9xZVMZPOqrcGn65+Y8GFtwOH4BoAgLBQqs7xDBDD5VstD2Y3NjUeJ9Z6Ql0oG9kIU0K643hAekB
4FooOX1Lu7R40zG1IwK967XcNy3ZhfdvxikF6pZT7FtI7v36uXf5ipOBPBUdEE0yHFuyKY/7l4Yo
NAAofhH0f3fMGVDk8O2wnJMkhtnR2WjB8050LtDDGgOuMd+fHNNVj7OOTlJysPioLAtafVbveDB/
Ht8LPId5A2Yxolh/1IUcdPjN5wxEwSRgFzsP5XF9LOJFy10flY8ZNYA6WMcVV/OQRt0Gx4aYGX6S
AV/JM+me3KIux3rf7nOFWZ5U9x6+IhYVHX+Gb3nWTWeQf7xbUcvIQ2yf++Me43ewCQjBKLfBAUYF
leWoGVR3mrCNzWRIS/HIFhI7xkhBVZHGnedsSdMRC8cjvPwx/59+6+bjXHsxXsHsuptauhNQiuiU
Iynm+IWhQ+GpfIqVQM5/K6hY5S4Yi/CA9UeBRJf/1U3NyirN/wFegTfqs9cwFvx73WfEJLZmtXs4
OJI1wr2inGzGmLlGkJEUGMWbKuYCd2XGPNzb2BNswAZZloG1jsIXyb9Vc32/DVs2rPiXkbgowhkh
EHzbGwFxApDj/eMg197ZCEm+dbokMUTCpHz6ZJ7ne1UsiJ+nYDE8oKNqLBxNhFoiKyMkAaNZc/LN
bNnGPbG4vj344wnowZMf6ILqjWnznLkn5luRvutgKeNKip/M14CxfpcDT3iWD/nXgjd5DrgCnzAr
GAlewBwXoLgtVIA5Lb8sQs3oTDOoDNMehBIRyXO2dRWFgivNPhhUWPikC+M1ZTgqI9dnLla49cqD
1SqZyE466KRgCzutQmi7+pErC8jLlL3G8sTivlDPXa9tBM7UlI2EBksxoXwweu5/yt521QNn/a7b
Peo2fQU7JnDofcYZo9jzeT3F5KSkzmgbKxC8+ArYhveEGsq91l3pURxf5PpttMDytA5IBcZ+4ClE
atCAcAJW1sYce+/N7yCz7Rz3l4E9BSxk2dOeGOnXB6Wjk/uSmiauzEsEw289r8C9o2Z0w7HtLe2T
r8cKYNxTwk5E7Ft7JiqrlwrpWyJM/zGp4r5eUGeNMFt5AXdE7iyLtkpHLR6FNyX+W+A74y1/tgoR
CbqhqMn1mNkXQe0R8w6O2Ubqi0TrUl6yswIcAoaGH3yNmF5oTpcUPYS+sJ+3jqgYYB8m212NK7bA
jRDMzvlgaPSOe+PCi/dbQOlN30fwRMdtOYyOYneIBXEvNqg7M1JIRzvj/5BcXIX/FFu161GWhJfN
Nix3J5IJmv60c9mrH8+EdGnTlj3qmvSd736IjIxrz3IBMsgKAXsryBeZ+FIvaFV4hp91ZQRnu9rm
xo6BTMp1pedwMnPSI8R83oynHfDmdG0Azc1foAAgHLkJdhvGPXirhTRr5fjMDBJTtSSDYPweWpuh
qISAjF+vMWewU8ccMsIKR7OFnco5k1iTwEG+DuCxu9c75iReX8EOC9dtv6EROPazjhejqpbOU1sc
r6dw9G/leUeMEtQLaw+ccGT03wnLjTzxZbm69WEOnMw3V4GW58btHFKczW3knwZDgcuLBfGBevfT
xUEvwV+FxnukkTKAadbanhKnzCfbTlBDKU0mAmvWF+zKXh/LCEszEAOPMlqoC2L9S7nhvElf+C9B
kx+V6yvKIsIPCmxoPSMPeBSoDEI1pAURg84umSpuLdHkTR8BbQSjeSKzQikhBQbZPsYgau0v6e2r
BpxreT7xC5MK74NihZL1NpxPSKRh3ud3hmyo7Vg67TLKyv809QzOAP7zYx65XGCrB/7Va+CRRt2t
60nklEZW0pd0vz/ul7V/o2fHxldb686K8xiYFoDlJr0z+S3+DMpJS+lSHqHWX7wklAuiBKswWmTB
Aq/V3Tsgk2WJFcJUh8i3v+1Mdj03qBStfvKKWyvJHQ876Lss5TIDjSK/OAm1U43ncKBoUywCLroh
qhcyHLstRwTQD9vDqj758l1wTuMHA6II9rZNNO19+uVm8MDXaN5jDlqAkLXUbjnxLQvBv7uFUetj
RuL3J4OGN2wDrxNH667C3WNtDrIz6/HvNTkKKa5HZ4RpRLtWe7NkjZKMHdR8HxZlcRerybKGuGOy
nLgf6EPU3YLrZN6gM3cHW2hyUCe7nlQHWahpZ5QJpli7KwyKmHN/j1bA5djl+yZ9TMASxpzWtJhL
JUAU4nIxD1Oa6m6u4w5U1S5rJqzNnxSzfTIE8Zf1jAJXcazey//WMekTmnnF/pEw3g9NN6jekraK
qardnYV67xMnaHp340GwRCRKmb5k+Szovi0SOpVW8VvCiI7icOga1mfeHWnx6ze3HpPOpz4K+sWd
0SkDD7i/20nfRMjERDQR392XKgKDPyy4LS8oyZN3Nkbz+77AXOnauaCix//Kq2blD3hLpOAPYcR6
Hqre+gUuuY+uaab5fjGBRxFvqAdQnAgxV3+1/aM2OujGC2CTD+4D68iaBoreRDDhHjd/O4F7wsG9
Z7es15ERX6iQSv36lAxdVLWcqR3JvFz6ur6fSJTxXpavrQTxwXXVjPNqrNpgZM6YgwR9xRzn9G7y
s8R8Cq9wLb370YitfYUF39r6wWEXzdCEyyVtK2Uhp+rPvKF7X+Sug1V7l9hNzCUYu0qpL9euvoI3
O2zWdZ1iL1Mgc6Tgv6MgYOVEgaNNL8U2RbBPpiQPulss5OPcAIPBUfpieTCERftJm0clJDfQm8Jw
spQhkkK97WvCHoQJowdGZnRcBbWhGlVikA1Kw2VGVFpRhf8t+SiCCt2xfnv4qfhZqLcjhylriod5
42bngFQLz+LVQoWdwyEEW4bKWssbiSflDfSc71HUmmfoIqwV6n6frmYfE2lwtgqHbwrp2K9ZnSgt
eTYMXbEk7HRMlnWAR6iyaXFaRkkjgQhkNKXNzxR0LxrgXrjJQndQnAYKIsuQ/oCq7tMoH2A4E94n
wPUjmwHeFG7V8/Tn+1YWl4bFW2smACNjSsn7eoGVxqRbicQaRfxfZcVCQs6YoB7AS38IuTavRFT9
kFbD6NwKrr93/lpEKxk5MjFxXQ8RaiG3E2JwAHCztbjQrT3vgoxQA1fYIO2XqFwczld/Z++zFAa6
qN0qeKjk8r0H4hC8p/Z5hOlGFgoU6/BjROJapjS+RSUkITPqZzPefbxZiRiWtq1/T4sAa44raZY5
aTHz1pWInpHn9fc04KcWEo8/rbLeooVPHj4oE+ulEr3JzkMRvLYTfKaCu2XNtf/KWBRoroWKuOob
ZYUgL+OCDWvVsq/Ctl3Ua5q2NzZdpghKUhnYbc/L74RIOrOWEmDQS8lQIi4zk8yjue3uUxbyoMd2
TPrHCdSayllXfd55GBxOJ3k86fR2WJz9V6njhNYHPJyk+rmygkEU6iHY8r0isTZ8vw9fg1JDgCl8
2hQDS7q6UCJKXku+T02bGQM27JBuN7ZNpGDIugfiuglN4DuVFxIE6McA83a1d3HlIVUGekoak9+u
+ZvL6MWRqjvkh2+WvYUUmz051p2aUvMGJUn2VikLjB0b4BaPuHJHxR5UyGd5mQV9yiaztWQ29sI+
S/1desHoSS10M6XWJKgmCTAbIpGGXMClLurm0dJ/mVWxHk9sQ9Phcw/mguJmwRrd0cNbsK4QC0mk
7v1y82Kgh48mvdV2crUT9hH7nX+dl87YUj7eWE2qfKlIJ/l4fi88FWTaKP2+CgN5se7+3XIuxCwK
4TlGpl7bkEoHpFdj+htKdPejiGTytnrP4g3FyVmJ8RVhOBLnkH7Lx+MadSJ9zi2aqbyAStImQXRC
Xn52xGdBXplAohRgqKg0SyolTrePzNlHbttKyAqvnB7BMKKaMIvmFyERTlECwJzvjN2r8YuZaSvS
mLpjuI3x8ag0GKsZOKDXcpvd0F9/CGA2+/53jHlS8QJCeHNF0k6UsgNW7kRb2hbsjLSFCXQMnzCo
gpv15aYmKJR+XstzU+KSC8WxX4/g5eMT4rnw13daZLa+wqSxmG+eGRigS2PVaFCnIP1TgUQ+d71L
5svnbT/AB9AMLMyJcsq0vU2Z8Y9iZL6iJed00KBvQ3rD/3r5WNKcF9weKtGnXYgWS3GEBZZcwLVH
VblPaUPC/SEwYD7bJP4qkA03kJl0KSpUNUm9GzdWXxBvrSz3Xrkuo2WLr83RFRlFtdTTSqsaU/tI
BuaWbWXAKZH/Zkw/RF8zaLNj48dNaA+jUhLKiq2cofsyty/ZSHN1jba/ucNQRDsOtCS/is7du8zM
LQjJoCNX3wPKUUwMQaXbzBTfakuBtQP91pz/qnpgmCarsaHZC5YJpRBs9LSORt2tgOS0UtE9X3zJ
z8VTw70M32JeEK+NRYK1F0CRjxkaxV7AX6AuakNd4yW5Tm7rworWMSXDWixZNa46lWAZq2PsDDkS
t32bGYjacFH25kIvtlM8zleBkLvCOXJ2L+yGbcIPCeAws6M98A7gE5xZnCckxkYxj1ujofgDxzGb
mWbgue6YRP0G86dTmoclHZDqiFvvrQQV2CtKSeETrsBEULzF2tT851SWwDai9cveirUg2yNbivFA
spuQ4GupXKtOGR8M21Z9QMLFRar/XTbw/PdYYBpjzVnBqs8nPNxf/YVXWOXg5Vxt3JhveDFculls
8+qCS4ghHTXKqKmM12q+f5jB2WE9qv4kk70SbQjHEdw7PAUe8Qnqp19tQTvUCV1qJm52yy6sgqQn
c0ZqIKoKBzpQAoKXw9dZnaoNinw/9LqInnb2TkOEStMj4ynJ8ZBRldBoI3W/B5v0gnX/n90XftbR
LdlX/px1Epz6uN0s0EgLXaiosfSWAlc2RVp+qovfDBUHTnFV0gvZcOC9FK5RWbUeaULcD9DG13XF
8pTTRzzP7V5QjvLZP2Ea5YNahaCQ0Ahqv0776YosVEyLT+K4EkCP9lzf65re9i95/s4j/3qTeztM
geEhQ0A68E7bmGb1Rm67zhjTt7y3Him9mQUmXZgRWvb5XXeTPaDaQ0YNTxLZDzCBl+OtpgiY85BO
/tF2KJQVdy4leUZum4gLuY+47GfbEfW+qZThpuNj/kgChaEz234DdelaBv7mqkPN+sIl9YqK3Zvx
oM+3b7HmOc6vEHkmqwGtqfJ4yijGEUPhumU+5zS/D04jnmNNDEEF6HpYJI5x9LWsMO1mWy3e8bPP
N+Ol0yhFg6DNM4nK/JdwiiG9Q4rPasBMATkEnwukRMPxXWQ8VU1y/gs1Q0jMH5KuTB8vwo4pBTKD
cpA3jrbH0H963xQz+5ArPpmXB9oga5x8DTP0N3A4SgkUsTHQdf/AV9TMRN6YSchjI4oo9n5fBr7q
p8Rj2OxP0yHD4kqvueduOP2/75m63GAC0ygmHEpTQkMaZ1MlDTtVSszddg4PRnpXgJmpbkH/4PO8
pP9qfmOjNNDTE+XSK+qRnEuct8RDrqYYPfuANyG0oY25bYb5lSn4gEO6Pa4xROV+JoTql+p+uHqm
HjKYfNN4fZL8me/9snq4WtlvlqLl+rj0EOtdZ2rT2bBZ9gl4lxsD+LzArggogCO+VD2jZK7GIj5B
jo/BYOUzvuJHABUR9+e3WtP+NnkB5DEdkCelPaeKUqfaXmcVumj6pBnJWlJi3OPOmPtBbWNNuJ/w
V27kTYVzJQQqGCKeCinfdEk/VXmbQxYgBU6ng67LzPoYw8jmYtgT71IJndqwZo1AUGBnOW61tdtt
/f1Jb1D1cQiJIzBlQWebhfM/iGHe2Vl+4ayIoeE5QepeRMHgLNPRqhz6oEI7WaRxtHqdZANWaxAn
kZOSWTnVeSGp7uYC6coMzkXb4GmDL9jxoJOc8JonXE/kFNzqtLptriQgWlN37seY+/tK06Br0kgJ
418UpQV77JbyXpE7oi3qok2LOiYhjzKU03y9OiveuAZlJY/hhKKP2If4tgGhHMtUHt33dym0OUFX
YON+vt2rT8jSVN4RvmwqUjJTCis3TMtIQTHr7Cbi9UWcDX/l9LV9TWQEbNpZkLQGUTR1DG3K3kkM
IqtoIdwDejuKI5XLSKCLIJJLTihYVVS4qKz4BDM2xUZoMsg0+l7x2NzaUJvkEol/oB29gzTNzKr0
Rp8gTFLLEk0ncyDNQ9peKxVDangzXACjLt83v5rqytZvw9vznO1FS6Tis4miTM/WfLKnYzg0baxb
8Fi6fbydJ+aiq5xwVYdaH3g91EUg7NAJqRXWrUeW7YfWhflEolJQovufcEVHCDuoogDzdd3Y17cL
OylRp1WoYHa5sALqbuySL+8SQ7AGljc2BmU8/rIeBX93oRx3rr+DLfIhyjUb5Z+yiEQmDbXS0N6Y
eQWDZdt/2YE2xGzkAMzfBNhD9DoevYjLUkJdti2mbPOmQYf0lDX800oRC+X9gu1g4o3oEFcLnGqm
qCy/BmSfip8xTOyxWP83Sw8kus0BPCXoOFTjXbcKoPsVTf4MNdlARSIcHZFnOcPIMotIcRgK6sOC
ysv1fRmfiI4ERD9w4MAgwjToIiFoAbNS8DgFzP/U0sbyYDgKkpOEYMf8hqibzSyoKaMDVDHeBrzO
Tz5QyDM6q1s9kolL6P7MqycHMlA4+U+TZOTKHdfqUgRUxDXvqsBP2Hz/HWElNq8nGylE7JlVGrFz
6TffWpGDMviO3jVv/I9RYS1cirYbRdxo1iRidPlY7BpCNfAcRLjZyaeBIDGrYtKQfBm2BEWMKxeO
6gxhw680BrHh7DwDKt2FVd/8FXZYaZuAERwdtpTmq2sbFcLFFDs41vafTM9QfLiPI5/iDyy8BDzd
z8qS4Kr6Wg9f0KPKX6wyG9MnCSV61AQgWyz4enmC5SyMwpGjtUJAgiqf4Ad9QxRLek2pjhH0zd3U
2Wb1xHyAJJDtuaoEyZ7FsN6XTuGlnkhQNIVxqCnhOtpUXKtcpGOiLD937jBI3owr4eVT4ofkkFY0
wCXfyY2B6yMD6hsX73tprhvQY66NgwpTKwcrBnRbp0cTcykb1DapD6aDMYqT5JmvZAmro9PH8BOL
2S3X2tvKjsJDWw68d9BF4YLNsHHtkjmzUyoHDG4SJS8LXugmHheuP7LUXKCaMp+Mr9tiJz1k53YJ
4jdYwZjmE4NbR+9Xip/f9p9hsuWo8WR+lSMJGfjcWtTqNfxpqZUINpSkmV0CqfwHrgWv5dZqBrC3
rXwSAQd2KXtacfGx+GPIHtMuj8/TPZG1sJLsA0/9JTiv9hNX1PDcRyEkhx8ZMvy/kru7coRamcsg
cqS0y1d/JAYP+DCM85AelOpoPNdEEuedDgJS/b7vhKL0X868XW3U7hsed9DewTPFp63HSyVJPc5Z
hfiGMjKFKJUlCbfYqWQzHPz9R37WJHySLIAuXkGoj1ICEsvBvShFM797n6RcFckrFHuBk7btyYPP
6aLjREBiUVe15X1DTl+MNPHb8/Z1fJFO2V8RkNlmTV/V0LF5vDr1epGNZRkmMLrSYCdTqSgOJXZ1
F20Z4LY/9OCmtJjiZ3tD1ImGMGjnqE4zPKYYzb4EnsETCAmo4e+86C3fVJI/TOHDekDTJJcKpRkb
dEktY+e7+9Fw/HSDVTw6MtcVwNcsOwX9OJHM74hLwUHk8jzs88d/gK2x3ZvYy1SwKybBNDuq9DTX
W7VB44Qwc6MxSfNRGIPa2qcqo31Jr8mRy5S9idEVMmdqOF34FmghC/QyYm9pmqDGf0VwW16iX9hu
3GtLlQmIZE5T0p/m6xIH9rNhtsZPK70Fi8u+jCFmjdVumpoXlF4xwHnufvUHzU7QKLGoyiyA8kjg
PbmjbENyLNthnSqQZzFr44DS1kU8d54vTjyaZSovaZeBJ88xaKPmCsHFd9WaC0bjG62/L9GrNRVC
pY5NuRIJSDMi7mYQ1+WFqURZ+TKmX6YeaEuwsrj5ELfDOitAMeTDCR6wTzRZm9uHlMPx0KtfsZzu
PcNn8AF/Gyz/irT2lhiAq6+6DzbORBr2lfI1ukWfVuNKI0PNKkfaOlXAFi50vzrO6hwlEL+JeSlU
L4adHLz+OyzEdM6L1NzFR9eMBqCyBE0MCV1ncm0EOMkiqWiP72H7hTYgQbf+1tnqRC/0qpxTffYV
Q5HtJrwgeL9UOQvF//ZM7kEGtkuguvTLdX0X71oQbaIspIanNR5hkn7Nvi6UCwxU9BDOFMJjojE3
2DJXRnjzTgynGlykxWyI2dkKSijg3TpF50ogpm0ejJi/+835tX1PZP82yJxUOvVYrDJV1GHSBtf+
TjwscctZUPTXNjsz1svGyVbhRcnJDG7uQCzBAIf3Db9CxPDLNMZ88HNnVUcRnQ+FL/XmTAVra6uy
ZK93vclaS/pO/2gj9YisxoiKeh41SyyiMyZFF1nHacUUNxX+goQdu/iWATy29B8zcQjYRmHk7wPH
OqeENIKvO84Fh0NjIrJ4hXlUOEXze9yoVcWMFY+VJRELmVZQlKoJOCgbksZwz9w+XGlLmuRbNxBP
VdPk/ZiXqJFW4Z6/vXcr5B3YGIL0kpQKq7lIf0NIQk0QZspNGUPFlGx6k20OkS7Blc5JuU3L5gAD
pfHU8/ZYlf3QfpOCDcf1OsAjXi4w+Slpy2+TPgSfoVZf7Wx6g1wxwFTS46Uez8AzP0lZg0HcySgG
3YDIRgrqoGxyaK9i4K3uUrZ0znFAmn7f/lP//w3rS3t1ODr7kuCOhfthr9EdoETpPPfvTxRIQBlR
vEaPO9uU4X4OVm2VNO6wObtPlfV6VBKaRHJjMQW3jZOIJi2bNL2f9zrPCtUGAg/V67v8yaJWQSP5
3Jk/XOjpak4eGVo45gZTKac7BM/6obQtIxLn/vjHMW/+umtH6ChHBHR1EE1DbBtYY5EgcjqvA6tU
4VLJexn89zREFQlk/F4zQ03RkKaDraRXlW67OLLx+8Y3kSMds4FSVtDHbcIk2cIgdx6IdfS8rwBZ
z6bNilD3Wam8J6kiidCrKphL86HUkMxlkzGom0qIBzhz1b3UB2XmBzeOgN1e5fxGxlUHoF+Jop7/
7dZx3VuiORhH4SPbGsbQ6Tk8qrVmpESpDoLEg/cnQhyVby6oO86VX+/YtvSoskJcoSrZgaQnHI/O
GBCFTJ3q4gkPo99VYEUwu/t0T7sp9BY6YmFtWVd1z+kpqh38f5WdyLnNN3jYoBlJHxB04H+ciMfZ
mAGxPVRZ+ccZ1TOiMJ3qdBnTnCqr9dRBStGbgToPeLCyQpSPwjQpYcKNjy6GRa7q+uOKCaThim/m
6Be/ZvjQqe4xKADCVMfDMB6DT7njC5dy24Q96irmY8/rx9e9Y77sMA5Cnhk+FRDe+Hqea26taXRM
MRFVWn5JNWvise37oBZjpve0TmOJPCmdVXyRuC1ML355fJjV0CSUhuVQnhQiCM9tibGOy8KboGMV
Q8XcO/qjeX99E/IrkrbfepMX6hNyMXKt8kppOmAm0gxAb+GtGLZUzmEXCFb1ofdNcfiKTazuMbQe
R4E0M1uwBsNPzUvHOqkR/tU+eVdXBn9k3tiUdIcrW1SISPvrgzZ+/9EuBRlubS3MlPluPhjmSzId
xTAa2wonCjiHi9yo6gFtDk0p51RLwsqZvqc5e4Pu++XQJpKPeik0EMWs+LgaRLZz0SdCtbo2ETrs
FwCMgVXumssPG60gvPx2mrpPwTBDaCCkyLCrov7D10Ug/Z7CA8uLNr2KIP/LUA3x8DbhDoNTsJGR
+FGO4+Ypycwu7ygaGbbY2q5W1q4CYRkfTvYFp8H6AvyoYsHLre/DKUZi7/TBQIZ954+OKlhJico8
Xt7C+W/yo2KlZOipEjoMjip6DnR7gYBCmU5GzPQi9XGPipj0QrN0PDzRmwt8jMKfe2AURsL3J8+A
S2XDR69yEz2n62r1SYYXtl3VMHdiTVWU+w3ovuC+e9qRo55B5ECQtzAEjWjVrFCCUGoLqJd0L6cX
DpL5KJsaj8Rn9sjei/Vobv8sME+uXE7BrrjuItXLMw19L++bqkhOFzsM1eheT1ZDtFiLJjF4335k
Z47EbdiG9fD6I6MxolH/4uIUrefaniSWe3g70/AW5AENmTg1jr/GywzxB96eXm3gCMHNjJ7rvPoM
ZqAVDLHofqpNI9dbZ6Pwb3m/AH427tmPxCiX2aAvYJ7t1lbFlLXgCFvvq90lX92WFLOsCpwzcfQy
e9A9m5ksVxRLbRrCj1zQCBimgZlDaLq0khU05GhMDIIaeudnVcN6RgKJ8VHUpCGHwUvuKizd62Oe
8JTyD50nujETHTwFjPq9lmjN+fdXUwYOFOzXGKxsMmA+fFeYBlxxU0cYCnv6IYJe59C+RHHzp4uh
fbVgl1Crz81eah6+3MedfUmd0maDdSKAb1QQ9TLyA4zjhLJfrho6aMvGb6XttTgIRxxBFTd5nyhq
B197ArpCw0Kb/wK4avyVC/fnMuMEL7sspMOXTK6W83LKPMnqzzhYYSgIfVKO3/03rIJ3k+pqhY8c
SHrF9vTK6N8qqvwZ5I/wHPQsxC2WqSW9QwLNj/HwSIMNt+d02ITlaUSFp+U1SOBtuAIOnvC/db19
vHJ4G6/LeNzZYO7QIYWT7ArLqmih+b0nAOpAR5sG75zUuTCu2DLIMvUEo2B7JO3fMY6WGhTlsdSU
LDE3FFRsiCqoAAIoRvZBivOYd7G8DIDgHu86telAwJRi2c8MesURgGP6RiU707tirhqyjncaKWpV
ZA54gYLM/ob6lgI9//Du2PpjbqLiJYhTHrR25OT7JCAqRv3yMBWvzt2e1DPsjHkvu2U5X48gyx6h
vN/n1KM8j+bW7G4lzqaGPGhMSCaozKHuNjJ0CSgXM82FCQ9snanxJZ5b26yyMQzjc6LL9cPYsUy1
Hu/+sIbdVkiOAQ5erhM1IrAnk2xi/JeyzAQZ4JbwZd7byuzGzPgmML95a5PZplrlrKiu2zxxca4E
fec1CrtrNHz8UAUX46N8LT1HjwjIhtFO+RAV/SUx6zyNSUhmoLN00aixXJ4sQXrZNKul52+BEcjD
hlJkd2A7uk8HyuL/5TN0MeqqxRwPt3xOrwLD90bD2WrHohrPExyuxnkiUJZ8pwlpxLw3lXQAJKf/
31UunplM6Ub5YDItXlimNEf90LT9dRLYlilqR1JGHKtn4gMik25T+pUNXQ1am1bhdKj7IlBm2O14
/GGFvdv3hxAGpWi8L+sBwPCL9+XnIb3rs54CynAsLC0U7bcBBnqDYEOLVrnl4LyIEzG1xIDzilCs
HOWEu7gUZKpofhBfjUBDYnE6S2fIOq/aTYaRmTmv5SawVimxsOeg59yt5T/FibX0Q8ZCuVZEekpF
Al6ha642gvF7Hf39FWhTIV44hW+X0/XEWaMHcXDC9a3fWD9ZqfmawARtHx4+zACXs4xUdzkGlNpG
BkddxaHuYepp9QaLMWbPCivwn6smTB797EjEea4iB9JakM8iBArOM+7m3jooPyYNum2dN5PS7y2Y
+fhS+ungogXVxZGNO3ZYqAuCxWMjo9XxTGePAVh6KM25IBA29za3X+LPt6nz7IOa6HTXYeLm8O27
aUAvJ9g2x55EgqkHE30vyk+DiUo2xJsP9xGPknhx5z4qI5podhNz00hTiQCKRDgTRC2Cm0M/OzUI
+FP319x7RKP0iVAnBv48peILmeA7V3pJ9OxHu5nJzWu2p4RJDLCJdZDIrY0VKeqwbE3k+lo9oSCV
Mh2iLowmP9M9NOBwcQPsKkanzXIf1f6br1YKt6OLUuaKM5WCIFhQUE/VZhF2hMgPRFXUr0jI3kzc
mrQq0ovfycJS+jAuOlhOmzwiZX4zPQT5tSPVHU0jx4Bf33uj/h9epKedBKQ7B7QpBhKwRdHNgkRL
xDS+HiLenufOZODGG/Pi8bxPF66GWfczvO+qtnQJ1bduddivuCp1XS60I0C8QGEpg4W2fLenHNTQ
9VV0tdtnMF98bmxfB6gKm3LDbNe1OzbRM5yUeu8F1+1BUuxHMZg49jwRwoFATPlzFqmPONLFZvA/
gsr6h9XayLJJhWwqDVegx/xrKkbUDEKRyVmfmbANauM5un28ILCUDu7UNREU8XrMQpWKv4ftotY4
+R9TPoDtI02aYMCm3HMynld9o4Dvi53W1Sgp5PA0UA0jX1YM3WBZgoVguNbJAsi28czHT0hf8yQx
I2pGlIVf7wM43CjeV2yveENKigUx/zTtL2iItUMxEbBFQJgUoqz9hJEP8UlgtfyctWmP7sjDyN+g
k1zTlWOVxfl5qwQTdmv5cKI32gWRpmfPz1CcZEl85uDxs7BqItuTiLHYUvF/Zg/Jm6AvhIX+U8nj
R7tysTsUziU2aFNrqx18BnboojJwmIdfJhpreOaf/Jc8lt09pvHINwCcLn0OUzAFaXSXpkR0CJxF
ureD0dWDZeBGv83OGNjv9HFZXptkUVfaXOHjk5B8n8n2eGtayMgz2ZFY1gr7PzuwbskglgrRFKfA
wfAqcN4KXwTQWoJYDP8FvRhunxom/nNSeGIlztsMb2fV61wboI9m/hhqC6b0w/nRgtF1cTEaYetR
Ait/EDGg7NIP0dPLevhWamtmkVhpX7V2mKDnTzbOdJSnQRJmdi0Jwbkm8kkbN+2JDUDHQLIhOncl
IqiY33zyzC4PslG3/CFE84lE64JBba2ZdVPZE0sQFeW04/w/ivrsheaKaUnSpT/Q8628O+49BRmE
UERb4vL0fEXoVxuzzxvARKSc42959SwuW0wSqLbptlRIbC5eMj9+JHMiil1NIJ+U7p+G9/98v4jC
YXsc2OZ79AQlCyeVwnjoO40nx+x5pR1n7A5JF+ZATETP8mZF9zP6hyA5sbnQYFztCO6/IJ+BH7ud
N33/8RUaHlfwB/SHDtA0gWAF9ysCj822DSTwk5ej/Urea2x0Rd2F3hfpw+WW8Lv5tSGOgkKiaTfa
ga/LUiF4BIxQuRdpNNoSPdBcex+TY5YEow7mUQ3g8tCE2h3oXiYyj4lSArGZfijvT4mVmsSCdfKD
wOi+2CGHswL8fODhHRSx9ZLJ4H1pybdYQ1PNy0E9Voa9j8q/zqmk24g1pWm9ZD8Iuug9jNcaun7k
j7bRLunFmJpGhMG0icFLJ5dGwuxQSbnRVyBRcThilWbVQc2r8kCStaw95Ck6vhLVaJg+Q+uaaRqX
2qzGDcZzVZm0RIpApevD0pVb+XeCvJ9eZ+daOziE96052aHXqBi0Zlzn8l01VC6f63GIGMyqaJMX
Q+ionbRi5aUbn3NKCBznkWofGTVJEL/pdE3pAUri8tK577e0284W93CY8hRN1syxhRfsS2Eb9e5R
6h/qrswhFw4eZkC1jGpEtzjO+UuBtsGomeSSSqD+FrSc6C4H59v15mK9cDDMB1g7I+Scwlq6mrAo
qpG0sOUBqEYbcqxT9D5ivQCBQxJkAqpyUQRfDixQH5Gz2dHAm3+tkHua2gc3q9sq2suIpL4vDmCR
6M96lYorp4sA5lwWM2EdQrXXEHSJxyCJWor84nAafcs/RStiI6dHF8PZgPvIxNRo300YkPhZrCkM
utpH7V3RZeBPat42i67YwEyjX53C04OwZGRPRr0LWfVRVXqAyU8OrXXyDdD2vwdOz47G2i842jAY
wt8gnffHNTTAkZtPLkS6FBq0alSEctQkK0hfU8SSZZc+NdNCFuCF9mVbCxW6EWEAslydANZjM+dT
59uDfton2U108tNJJuSsSi1NHyrgee9axSFN1IxF5t+oYiviST0hUAzsWg4mMktbS3b1cVqx6p3f
Jq2XDr0bXi0jwTb8VeGFYMxdtODetFz/fgNpeof2jG/P8asrqC1TnDkE83iSfotx9uqaDaMessO+
xsDfAyda14cazR2q2JWiEA6O5IQ+/SzgkvMnYCQ51jSuBdCnfvyW4qojI6hBRhh1uDcym2z2Fbp9
sgVbk1TBQjvVnRQ/yM5glqAoii2hpCpCY4Sm7DQhNNL6WgZmda5u9xVBziUTEVj1ftiZKtPKYu53
eOtzWBzekh5DwPvJ09wRiPG9ypKUBybgsEz4AiovW6Rg1t0+7oHkFqwtuMsEX3NeVFDBprB9oOTk
pVx02RHHSKttcXdtzNZTk8wGuJtEPMNZRMH9qMywdA5RYhowDMdZeEa48+9CQB8ddMj+OD1xbLcK
jWZuzGbA4BBje5s/B5hxQAqcnokXl6vMshK0i4g7YrRBAEhZwJxCxq8Z7cOupbHk9TnxdMk2BKHk
snu6eXn3vyW5IgQQEfVPiVR+Z4nY2KbNm4IVpAcUNBj3/sHVkEQHn3kcSBmGxp1MoD9jsztRZ3SF
Gl3fP39CY2Zm1DbLONAehnecxVqgzmImJhVBkia9sQHN8MS8oKGv0/fbwySvqdirnqiXkaLSoNoS
OUwZdq8yiu+HarMjlQVhMNw08xUYWo+NCycFyD7oOl9d2+ny1rwbjak2ru/52o8OwcSOlMcBjOYm
OegvSkK5oFze0PMY2U8wOsNN6qp5hq/MmyBekcMi6dK4nHN3I10AtP3/QRy58v+ZsbcSsTfMMvmn
nnfe/BWs1E5H60Uzrm84SCwc2rkJx4+CqNZYdyYDFzLcXxb1x1MyDLgqbTnMFqj0GSjYlmI+1aBh
zHNOM4zt7P0hLypTHsvVzul24G65zcFbBz/JNZdpiKHhs3p1AZcx8aOvTgn5caWGAKmOxC2FAfJE
EjsrBzTUXiNnhy5QXbRyg5a6Zi2s5dMDEUneI1HibB0TA0w4c6IAaGeWXSxvMBXfyjb4zD3gv00d
dhNg9tdxzDZ6yMEk1ZWsizD2f5yusxCJIO76I6OTHvFN2mykKSXFwZygrhLLPsVu4Bo/mUR8hSpo
KGmfO5SBp+PFvOWVk6hD62acKdJ1C8t2So+ZXvIh4kb5820+9nTLE9OoMRjcQ2nTV1JVjXZkjnbg
Lydjh3a0NKlOguBniYcM/Ue1NTEvBWcxt47S6z64F+yVMdCjPImmx5cXHp178YxaUMg+fnF2mbWk
X2ykJSGYc1rjjvHbFucZBKZxHYpnRVmetYv7qx+rP00GZR3/E4IFyO4wMTxlB5U8iqAiSiLpzMtf
v+/iy9we06PavDTXJX8lfLYN0VI5RAZiN4BmL75sObBtGqB6woYOdhTMDIQX0w/DBIw4tTHQ9kkk
l38il/txPhmMbP7FfY/che4iVAEck3CZSirzNvJUDWEyYnj5MN3WvGyA4DAhbq6PQ5DlhDmfIrI5
5MD2wBQG1lLgFH5PktLndsrjpsBpvT4OnnVZV+LHgpoe5gD9+n3N2Fy9C/Prk1tuChetuck8tuIe
ozKWc4n1mJ1vdi/a9DLpQxyAiybuc19YNmVh7Whmpui+SJDXFQLTKsrEAzxM1XnNeQp4XzksuJqg
jBvwtXlXvjaAGaiHfb30IvUFTUlDywtvRyOjR/n1sLsynFKF3wNwh3cMPj2kU1bHLIhtOVKK8sbu
GC+YuM83tXv2C/7XI0XPLT5F92Ft/1q7o4dgINFAEpRco8gXZSt/7dcwvfxBfyQVtxUd1KZqM9aY
jUPaVDQAjxhto0CRrgNf9Gj4mqeu8XrUQ+zvsMAgTL3cgL6fU1ZB5HWTSYPaZRKIk7ZM1Z2D8q8j
2LkrFOOD/xy/zKY6w2G6aZczt2ysQLLHIxnUT7FWEPeRMYWXKvSIVfd7mvraD9CXbbKdnzJCNluD
bJRdlv1uI+M/b6GkbBPCEGEog6hkeJtL+McJvscyZn0L7JOQWZpzj2ZIbgSvPEuviNalj0SQAsZV
5PIeh2DZdEdXPlA9WVDHp6QFPl166tIt04zVvRjD4a4b+qrarN3tH9TXdof7MoOyC4wxQm8yn6RO
VA7vFUjNtFS8X3X/NVUHYhrQC6izjY35ek3kt28n35MZRGsNJQi5OeVBPCnoVAFKm/QpVMuaX4rt
1QhzBy+HK921wLhLY+EzNMpn/obvdwCP0OugewFCd10pqiLUS6yQBJRLTwqlf6qOCXbXEheeK8Du
krZ1Ys8H3Cr3IyPSeQf4bEuZjfNlo3Jhv6y2as7nOSoNhE4eFe6x3eCOkuBLqYWElRheK1W0aDPQ
sEQu+gXxMJwpUKkMau79fjUkMr+5fuRdzAcyyMI9eBoPfmC8kdJfedER/TC7ClAPGrOrsFjoym/z
NoIOrb2nJUK6WZY5QXrqJQkl8zYwp4Ty0avdxVCNRwC4iCtaqJ5z4W3FOLjwuw/EOjFL04rovVvQ
mbAN3n28HBxGPndl9d+6eh6+lddH/xoqwD54zUJrSNn/y6O/QBBb/Aqc1Rquv7vfPhoGP37RqzDZ
lI5bF5LIpvLlM/FHaXCK2dZiIecFKRCnOmW8ItmABIhfW9jVkZR5hLBkQcUdXOH3DoSLnodo+e0j
r8hQK0iyBQL1u8d6LmhFWxK+Beo28uz54RksiU1yY56388rGGA6F3LF/JYu94GYgiXEH/PjfNAgQ
iqzhB34uBB13HRnKsgdrc5tIut2OYLdhzlCrRm5OP793N4QSpcpjAZZhG1WivpmvPVoKlrAGQry5
utUgHvs3WuNY0QzTbPnWSX9Z1nNLzFdncgtHdrBeh16U9cggZ70XEiMS+flTdGgDDN1gkZYF6Ia/
vTchArIyRfA7hPJzVB5G9vgv3sizI1CZ3M3DYsXAYLvMYuTVulHCfXi3czDeyPeIF90RoRie92Z2
KsDT7a3JQfZNE1CU9w/wGVpPinXSxmwR84pinVV+dgub2H73t9pvUekOgUI4qvK69HhctFk4lIp6
9Kxv+c+o44mbFd4/fCTEeu9vQWD7WY0XhlToVW0w1nzmoi1/rN8fCWS6Ng6zrm00UpMLxaGvGQpG
TK30KzosPDEap0fczJskCzkGuNE+xmsVux2XVibJtY5qQ5qGIeRPYvfhJug5hV2wn8aMOyRdpJvb
5fIvbNyTM1KusTbufYKhnojMO8t5PTFmr9f0g+BfwWwA5pcPeldjWbuxNWyr6pdOh6pJWavG440P
p75rwXNfp2i9HuJe+yxaz+OjVozZhA8UN3b0VXgXdKUonvRFG7CbiJhqEPBzTMGw0jlCS2E/8+Nv
rQwN9xMSW0s/bRjhGY25aYJbIKt8xpPihcf7OW2bL7moW3lXKa+ojBT2vfnW5M3Q/OppzjHpPrq7
bZK6K7ZJSRHMrv59RbXw6FZ2c5QJ64sQco6kdfDPfrvpI09zalQchCvA8f0iExUjhOrpU+T1jLBA
1Ael5boCJPxLXe05elOylFLR2ag5eAk5dtVd86wkqGCATqG+rN5t+SsXEwojOYswWqjiOA5mP9DS
AO+8q/Ltu7QpZzo/nrNZyPxsdFBdNn99lYJAptwSXwTKo4TrYzb1cr2mBUdgDesU7Dcz30NEzFqg
s4OwADbtHjo/rJmp+9Ww3LTiQ/IABpt8G4ka+ycJGDu10d152Nh3PNgESxpboE2L4hN6OoK0veS1
d/7Ww4sj6vcFyxAxd70CK1bXC1nZWVrvUG+dl6qUzHuzN3F2uTMPrc9bHjsD/T2Tetste85Vdso7
2ND63TEh7IwwL3MjHvsVmpcnCv39czWT7wWOlUZiTVBqxUhXnfWpNfAkuNeWI5kY9fYi1pWq4pEl
3crf7FcB7dsw3diwYv4dB3wN4cL1qBJSAALMZyiIOVVzfPytJjYAuDHzd2/ZJZqA9Kac7Q9OFQkQ
M9hansylbK594AhuXe5sD3VkBL8l/aKO9a7fAhoAlhP1zntWYwTEw6hw5EJCuNgnb4vYhLI6UOuT
T3nYRsWzvA64Q3nPp3C1KKbY1t0U0rQOUg2nyaMZtO43Bk12oxrcmkHiFQagjhqlJobLDHRjzPa+
u14apwN+i7zfXd+pbN1aXhK8hEjlhokbRZyZpe2/n0LVLhhb6FS90Czdfin6yz5pETxMWg8DB6Cn
oSHdt9DC/gHngNYOVWQyO/dp6tOTCM34/6dPQI2k5EmoZmH/VJ+nj1G5FU1eXRfe7c3zBfU9N/MX
vutyAd15mEiJtwcnJIrrCgrUP8lPLImIlW+dttKN+xNmtAmviy87LVA1sUiIWTe6+H0w5UwHPCAt
zj5mQloKA8DSYClzk4LMbYhMnz4QAmYA1uznxWUaGsSTone3ln1twoYGaxpUJx9o2hkut4+bsAfW
PQSJOmlJ76vKF1CHaBuHXP6NeIPoAzgT267+p9HLdF04E8uxhoUac5J2njFNnkvd1mVILstLLz8C
G59QeRJLCl3bm/n8P86/wyE0sI/kq8PUvIEKZBAWFsxcZHkspzNQLtxS0KwzQ6wnxKfDd0+gFSZp
kl2Hgdo1JehI7c/lw/OMbsIW+YfoTVJJEoQQPdNuBMlcPfnK+RBQXhfFtpIH1gIhyQ7de590/soM
CWCik2K9xB20vNmiORr9VcU/QtLbjWd+tFS10c0viv6F2U9j1QVX8ZcBMe5HQqjEhUV3oFbfYy4C
JE/N2G2azIkpdH61pzx+MH1vkhj7YX5HuB+BDTfmzO1tvbxEICwvFK9bZ5L+v8IJcEn80jitxJ/M
0QwiPC4iHejy2u2UPAs0VEOuJFisXD0WR18NuJDW9k3IDC9OUXtG+WfKPY9R0iHiETWQLGvlUXBs
+3cLPM4V/NXDeQLIPJ57DPM+orvhbQgONx4iT5mG9vMpyiADMv2Pgr/kOnNn3bCNESSMfSeke5zZ
o9M3g5CmUYErU8SACu6pkRngznf8NLLL4bebiNtjDOa0NFYyaxhL5VnEf/QaJ1RYsvF3x6R6/YA7
y4tIBJXjzzvJZtPhGUiENQDGex/SCZ8p0kOq2hwPdmqc6TyO3teHo5h9Fs98mihp3tbe5744DaBt
lFGXqburxp5jNcyK8omdQcCBoIgf3kntbFzTRXfgvW60k8//YvhWoSQHDlUjauDuZTAx4Wp2hqcR
MA6o7oXJowQ9E80zSf6RcksgypoCzX380Rtej3ihJ2fjUWETyRMuvtNouQbM/NAT3cEK72BABKdy
5QLwKFC6uV1JYgd4I/tv/UAGwW51bYwpzbsR7mkfi8CbsXjILLdL2E1CpfW7sfYfN3awh+x18b44
YfMAzpRn4tS3F5duitfftZXjifC/NiYZikXEP3ulrZEEro3xsNiJOqE5gkBqNymfxIlsmskNd97Z
4ZDBonpSvWYGvhTevsIX1z8Glvy3V4iQvjB9OWgyi4P87ERumUxlA6IjDq1hopBoM7vYgVZu1zRl
i2iCJ1k2MxUKyx+DP40ICyo+OQPGZ8AzlRoczVWNxdx83mkmoknR01Za/0Ic7JtFXbBq87dbD9Bu
KZKcxGDLNOTVp4mz/e4LYCiWBw/md4EygaQ+ZDcRz7zzGdaGmqDVhrk01NTq5uG1tzCjukOf0h3i
/aYqrZ90zQQ3kxLQ+PaNhcYV4OglbAJjssvkRpeXUpHALZaZsXU4LihL0Fih56hzcVz+FodQgUTW
R6Q6GiOnIhol+2ddOpxOdgU1ts9xSsaZPaPSRROdLdpf7g6OETKUwbcG3hViqzb1UNdxGXz2LCFv
5IGvGIt6xTCTo6gwhAf21Lv3DFySLCO0KIbu4uuIbVjF2OkMlgY7VKZfq4CwjO4ijRbxYo+/2NSh
elsgVzcznm+OVBzEn6mYmrx+PCrTZV+y8ponrLzE7of7hbeDmqMMrVNQlurt+VbnfvdAgzwP+2CM
1lMAH32m129lvPF5GEEdxLlz4BWjQRWb4jpeQrZHqplltgbvChUHDQaBgRLPB4omCiOgWcAd+i1S
+NucqojlCQWxvryROIz6CP6R7DTBq1NKAI0DKMOGuPC0QxOwE9I/5tZE6wNH641sfYde3QwUvZ7b
OuZw9b1gHmiFJFX1HWIHpkGDXEB1nuVHZPVOjDfV8565GIDFQCq3qMTaMyIbsIW2wqLmDEWZESPT
0XBpPuWeQ+gGWWtekPUblutBBJ2/RL8nJvV7eh7IFd4s8JgPgfvSyHZ19gW8fjKwXKvVS1jGQ4Cn
Y5o6OKRUeuwQCwXu9R+mKx0HVWcqfRnzfYkkyYe/b/muPZJ/zOdQp7BhwyVl3Kt7NhCYYkfJipVL
pXKwuTgbK79sQxO6e5jFTh8iOgGT9d332wV/OkTRptvWYaNhwnDfjF7k2lgGcT+19wM4r/rTG0FM
OVTUOPooD43pHp5Op5jZfTXuzON/d9kzVs39NRqof7wcwcHDQotjIJvvX0t1QNHeweCQsf6HRCjH
AS5pkKDEgtD2NUUqqzO3KrL55V2doy4uq0U381g8zVVgaSJ/XovIAlEhCD8Yl2RZvs+zMa0OeOoF
+JGmBOoU/SbnR9wFwRgMoWzuLN0l6kWd3DScYf+ZxNq5FVKwcOJ/3pWw1noD8CuyL1Ol97zudIhs
wDAiuf05ApRFAmWa86gj+kI+e/w5e+zzORLnGKRinR+Ta08H622Q3TSMDrJJ9GfT/xxSgaR2j1pn
RWAwvGaxePAedVBSlEU2lhwEgvCk8PxxTo6WZKn0mcqahJKk9gD2RPd0OiSsz5WjVGYkPUrDLoXq
Pj8x6Cm+Uk/l3i6lfxGCv3bqg1jI7JVlP7ZaGAwPkHNIdGOMyQ5alTPkX6db9//e+v58KJeFJsTh
bGNdzOqL8e12SJwvnV4FUUDWCx+yJxype79kx3FSQoWYkqZgUXXZudg4rDcaxbowNGqQxSBRVMzz
EYtn3vreG6P8Uc7qhUwlxs4pJdvKIoeuTWIEhTR4ljRbZSPoiizS76YUsiOxerpP70pGcvsCb2dP
ujcu9E3+ALHc1jq/B6HSpSVg4FotNYN9dxGcbI4Tc92XCiIRnmM5DwY9IQ59nvV/dyRbQ89UNj8a
sSaBPORRfvyR46T3sqTZUtUUqudD9nwNicKm4T1Zu7LdQAAu/L8H8W07to0hqTKySkr1JnmTgL8o
ZGBnibMqCAMf+TjBJf3CeB9ICR6b4wCFSSsLSo6HQUbHA0q2+zNhg0ylEGy+lU3GxGfzbfEhhAEm
5yINpuSe+cK6SrGlBTu/MD/xOJfy74xuOzEjzoph1ULaijuhgLTR7XsIn3tH0EbICw8Ky7B3P6l5
6c8TBKjkZZBKS9CPOHQvHc1gGCn2XPIBt7qLYMk1p7JdYQIGvLOxjHN1PSdZaxmmTCG05BdAu2ix
SvYKxSwls3mmvbizEJOZrzDTpVz2FQo7nAkBtdIDmYuh9pURh4R9zgGDvNNsL3nBYtaU/JF9JN78
3RM2ktQt3pWxq00k0urFay9W0RLD1clXgcE7HPveGHxTBHBEFCAFPcjZo9K8cFiXB0Dk/IHcFWaP
qURTjxTV2oYV1E0iH3roBS8EcVpjrNegyTwl9LYVXJ3L/O1Qwnw5Kqhps5FtWFQtxP/mG8FNFf2i
w4EPdRW5udgrLzyfW5SL4y81CeceC1rDAvl51I61zXEXPulXX6WWtqy5+89MJPWMcBqLHIi8zWMb
1uqR2Z7B6OBK+EXPVbVv8jzgF2k+xiY36+741VHiX8podsPBwF92/DpVVc0sCNNf/FFKG1IiyRe/
MXxyCIsMOfAPgfxJvsS837qlGjWln5lcPG7kUhQEH8E2YiQB6kE9rhBW3CXVMCuI5nc1fwtmVfxw
HCQ/8mDaK2yGo6He8ze54h8LqEz2dExSF0/bGeAtvgYDWffltEinANFWZjB5gHIOBLgDPgQ64P7H
a6qN8qf+WcqtX1PpU5+gdys+GhY0zrcn/eCbacMGTsWEhqW4UhDimnpn9vAVxdmXSWpA7EFjK5Tl
V6x/8Wxsc7F625R2WlUmLgrfYKNnkGitetv0Zbi2HWh++LiGvd0+0UcYJHxCesm5lVNYIEDvAL2Q
SvwLl0k5UyiVjOQxkj/LKbGzAZqkC/c8y6MHbOJmHatYjCIbZ0iyeuB+kVDaifGIQJE6XlYKVfEv
C9mlt3g0X0azY+90DFpK5VZ3KNSFMvzidk7LhKAfcfM7D2AiBjKPHieW+9o7GkPL915uVjPg2Wc0
CFc0s3x8+qHsnjtJIu/s+Wh6KSsOMZtp4n2PioD/vnRRGfFEk5FZka1Zzk/eS9w7FJBfu47AfFJO
fKr8EFT5n+FZDYfr7+udbfJLlqnPmIz5Ndu+0mD2Y/PnIDgVWNhLVRSZ2gw8+ocpgXIcL2FOx041
MW8F+3IfkcXDL5PP54c5qsHeNIGlcuCtoqDSnlAkC9b1iho9ZcbDe1hxXUd6UxJ7fPjHUSsmHPAA
dcu2xQukjGnlYuCJbHkTm0Bo61WfWLKx5j/xdvndKPuIUepjqdoqZ+/vHxIA7BIKUsWXJHALgaPB
lXxvF1VeCZaaGuoXKUnB56vyinu8kqHPIEQzbVwhEhTfhv8h1r0aWlXRkSo/OQIofSMDXa41QWvk
+5pwLtJ2uDwdmU56GEE86wybgxM41rtCZ4KeXgKw0RcH0BoGek+ZyX4kupztO5+5LsRUGetRmAah
uTR972ver/PgCwH1y+1N8WRfQRx1Ck0rfHtBpS3iRfhmytbrCzD15vkhOms1+f2r1MBEcQMRUPPj
MT0AhVBfRrKNS3wrbczU0zAg5gfzuclTJcbtPHz4r1lJUXguqSbuFmfAeLSz4pgGw8pfu7QvllvF
3sZ2YJyUshg/gaDTL9YfSe7yNmY1kiUs+eEfEJFVTAzB9CYfQ/uXicUfG15YwXQxdg8H2IzxmKUa
U5jtCXem8IEGjc7n3kBIw3huj3oHaXqZLI8vlz8u9TDyZXMJ0en7kat4GP0cus1L9XsAuRdEvnh4
259sVw42WnFsvQARtasHolrINkyMUjFBLGtXk50/dP80o/LqinQ/oDqpnIPGunuPLJGuukuthOvr
gGfrQYlvmtIRUhM9j5z3RgW7pAPNsCOlIUTBhbaa5A/9yRG0eq8ZXDThuGp5+5CSyl8lX7SGpDhv
dkNIIsUG2Jur/1l3by3jyTxEVSr22o71PbzlCiSB8LVrZePDItddKAwanvJQip3OVF0deblF4ONC
20HhD4qsne9+WQlhznEw605JrvL/n1MySAGxgJq2PlNPLTV81tLn4FsUfDZMUBARYhuVTsY2fzJJ
Kq1iYv0IKlYuo7sprKw3a8h/8/dLMv9LEw2rxh7z46myvn1Qb4p0N72VPF+eCknEtRFNkRq6JeTE
K0/JMoSd5UO8ABay9bFoeCfVyrwJWeV8Ni2Rj9i6WnpBRTLFi+w9MC+zRG6m32zj9BS7/W1XxUP8
C/sC9dLrcXjYjGU9165gPkmRsc5L30L04LnrYR1DT3JWksNnSjmEyOs4S5WMlKnPS/K/w61DVlx4
XljHPKIRB4CTHSejIMq8eCyD11CwUHBgH03GFcEiM7UefpNwUZZAXz6CxwNBExx1VMN2nrQfuuQO
AHimolj0kff5SAjwp1NLWOkbMiEdHphRr7IDIAn8Onn+3mYeQfrU/2u6mNEg8Q1DFAt4arKPipfl
kAuvtqZ7fVqLvFmAV2cNKWbzeynPHlONVuhSQeLs8KmresAL7BtyndEec1qW5hvtO7CdbEBkmI7z
XYMPFc4kghWOaP3bOo5Wjc8AfzCgKBeEPiutyQ82AaPpDZDI3uQ3CdnuYN2w6fT/uD8Qvq2FPmcq
NTuvHmPIlZa158JuIyIKImaEL7d5Y49Lk3xzbNqN2rrfEOJy8XhXnp1ERg/odMkR8v4hSZbk98xr
b8n4Tt/4iXPFIgtyFYvFqXmtSRj+H+gE89JI+myh/ZHGaFUoggwTScG693XpGqjvvWk8qxapwu0o
son4U+LQfgfQONaNlrovGO0N7NVgcvyCRGyr9nYJPeJ1sxm1zcEn+Y9yvo9VWDSBqfAGgeq4klAf
Gl1z0JlX7ZvRBHPP1yHWX5lZb1/0g+gvgaVVB1H/1RIpSCV5NzMn7y5t0+OsiZexuyL0WXZqgq7Q
OFA6OawZleVidEfee9dlw3d610dHRNbAEEBLxLwKZZ9/7i2mLuy1u1u4cse/4fQ26gZVmAPuzPMU
SR+jPwAlOKc2oFE6gLhywfVfP0zoRpAXkwDUI+tqBt8aU7aCiHJ8QWejF2AEhHll38iK7cpSE+rE
XvdKmoRsct/wIkAc5m41eS5Rm0cUCNExqfEMFRd6klcsCRPzZgIB4SBb1PjWYxig1OGMAd3vOf3z
HnFBaCcVdQOywh0mQMsIKJpRHwCY0j6qWgBMmGzPfE3fZQA66h74DvgpcwYcg912lkE3iNo9ma8A
8ENqj4sjD58F6AkNY/KiEcpT0i9gATccMz67c6OvXqfdmWi/pFcZIR2DhKO4jw0E9ZbdxK2TtKkE
YXMw/Qe+LjJSrXR9HofKdjxRH4Cqws/2IqmCdX/EJeFt0BKyco+O8mWstCa1TlZ+Y3tiysNHAUBx
NYhomuTpY0IVEsub716ypf9V9i4QbDrbGnLoXeLhWVlohH6J8bURVcwaQgPOlwIhH5aIb469k5t+
rgesJ2gqFsC6+J5YJ4EblLKOpEatgS3VAqTsnElDwgbUR4XrWMxVZGmTQiku0QW2z98f0doMizdg
5RgVMexet5AgwK+3k+j7xdA5pJOwPMehoD3O8YxfL1WJEeYullbs5XYtqUA7dP10kK8vG5WsosuS
293XT/xlaG7D5FubGNXYpGbQ6e5xW4lJOuUFfCAVN9jyBTyZzAURK4rCyIbHZtLGvxmqLpMhorso
oi/9vxiAeybJ2HSHjQIBTJOtWhSJz+QTL2hVKrcaxua//5ESvHRmC7h5EzEvsDwUjMkhfOa9/UZh
8AhOjRLL7Urmh5PBykGLtFAXM6/3agNMem/DL5ciiqys/s4Ti+IgRJ6DbsyW/PNyDEPYrEUf2vy/
96pfQR1X46eu67KZcYNREQna2ytZcidOXqvAN+yn5eQSyn80QTnJ9MbK795uvP1Ze22WbxpKMLEd
P2B7awkU6NKy56cW6R7cBlqWn1BIgqswSRP4RrWhvRT7iAtfAXyWpHiZVXRBCk0DYSGhYRLkAIq9
yfwUKCOJh2FIFSEt+1TxG9raPn/Dibf/0L1vQBfaBCAQSPVD7cZnju3DoCeBRwi8AUc2eH91yo/E
yXVZU62HwEkkFIgf/yxqT+TISRvRLbd1BUMieAtgmNctKVFr9Bl72cEdaKQJU7cwKiVtPqglQuyx
gemTMVs7TjS+Yqx+IJ/J94LAmBZ0eYi1bL1zTQyFAd5Z2Q6mmoH2JV10vhVV8HgeuuoTdYfDQL1d
/VZPehc7rJVdk4qMWNNllF6xLu7VBHT89VgANJdgTdmGibe0slMJf3jLP5eRW4F8EgQnOJjNx5an
u8MfUerjYk3CMXc091itpL8OViqgznuQEsFzhjpy9OLNDUMmII6+ftBq952rjzdktWI4DEuIkhVD
cXeXdwLPxUZNPis6jkSn4DvGBRcVPozK8qGDPFNDl7fEDfQS3YTr3sqr5S48CC2J2+0MBY9b8aNi
13LhVNJMtpfx1S5jMk2OIw6OeB+wJ8WHNuOPpyMQjt/0z58fTYcWZL7cg0VPbcf1UVL8ukmzTu1E
ctPU01UpttSSE5LISkVRqe/O+b4CVnswEuapnhKx4OkMoUvbJSR9tCfw8xwcSkSV7h1Ba3UpADuz
F2oy7HTJ7yD3NUmnZtm/9ssX05xrZyVKpUeO7wHai5UubTA3X7EBBYArjBj53gwiJBAP36A2FqZ3
YrWrg7TyISXCagyIu+wGwChQbOOV2bYfiCrgLjDuZYX1OWYjwyeEbTjRZkZrKSImPbN1z6cSv5VI
0uhmsyGLpKXkoHXnwzS6rhgtI0Zz6MIOTfy0QHKr5bS/Fc/KueJriyyeQa/VyqcFTNeSotQOjG8+
aI1Jk12PA1mD8gg5Op2GNQb/dcxTfI/8D0XjR/90kwpfDQUNslNutA1VlqUf3tPWfhLBSVaDX1rB
e2UTyklJZ/uwXTmwcPdNXqsZrY/ZI/QWSxi3AH2zn0ThYV/Jv+HDDkluXUOnuWtn/N3M4J2/3K+I
QTHmlKTiy3ZkB7jho58T1qoO8Nf7xqyKtEbIFFk2NSadAxDTJslddULOxBcdpUgGNK4W7nVzeyT2
SFCpD29uI35SE5kqhAo6TY8627cmKAnYJAMU95l9pWYDRqUrOgxoy9B11PUMMkHRyfpIKT1lErDU
EbUm4CbrHKYaGLrzVH9/xIXVMsW5bHOnD32YuXAwFcL43x1NQUBhHmHbg1Nt44fKbRJDBjL4U4Bi
4F7wVgrM2V1gACFsNXfIR2TI7illOFoATwS1M3aSFyLIkQ5fYDgfcO8GlXcdC2YzmY3ZuKmGx3Ur
xoZ28gtDYnBPmwxg+/NdT/d95GHdEgc0Dn4hMUlymS51aRz58QEjZumyZBpnPsDRfQDgNcYd4LPd
pcJvmsGuHiKaQwFmX3ZvLoQDawYz+JGUjhJ0ykzxtDJiSMILSVXuOvWl2ScQB2LtmtQMzpiEWAoF
cJdwaBqM7UPrlqKDpx3vJjRbMXidMOhOPxLPuB0zRDejgEhm54/tbG5f4TqLXa4M7tgRfRW48B7O
J4Zx/uzn11xeByjz1JJVQFn2Pxtpl02HXwrH6RDXNK4j8N0ZMcob0J3o5Fd2hEDicGZ16e3DALc/
0ZEyBf8m60XS2yh63a6Lz45YCw6bK8Q4JYynNqu1if/wc/Rt0cvjgaLkCY83LVAPYI5bmyv5YZfe
iCF329HD5S4ql4kntJU54bPEEr2OPEPmPM/AQ2soIRWk99POR6C1GtwvLl3Ij3urdbvZO+C1Qwk9
gV0sxbGkbGYHbNscD5NIag2lGZyXCmHctZQxppRHLMZh10pmuRtCnS1k7cPoauy2W8lIbYsUADUH
WLh2VIBDxACE7x2iysq44x1zHUcMxaOStrqGu5JzJGpQ3Bc08HIII8Bc1nKUIQgRatg+vts2SF8Z
NqQOnlkEV64dr5uZKja7ebG/w+RvTSdXNZmA/fgn5ZPmL9YOtmWODPttgDq6WNjwqLzW5aaqNMTx
rFxLUKJx2GSeFkJAiY5INe+jDPSykQjhyqPfnkHiuj5xSAGgzORGT0J3mcsSM2WxWmDmWtYIj3Td
UuOcYaUec7I/PSKUUfwFtQWAV39aN2lXIVTMMwX50gBds3tWgx14/AKOcwY71/26xpVyAxWRCsM0
3Wo3w7jq2IuKvTkkM5UH+tzPqcp5OATjxQojW345THGSbaVI6mbrauqX2ZdNE8/lNB35YiqsoYhs
vtFp2EpcGLka6f7ld9ml5FJnAsBG0ZCmU0LOOvMHwndPQQZE8qEInxYTstnQf9PGmJIytAGA4J4r
Hd6WHqGj3Ia8+5tzOrX+94VQKpqVHvLCg/NO2nsbMqsc6jPNBfwBNjoquMGsp36tLs8E6H8VP36B
WJDj/evz7cEvJQuJqNGzu+OXNn2UK8um0poi78TCJtXBnqgX1Q8KtZ4NV+9Mjg/AIL0S8y5But8E
PNsPoyEdFfHxUlGQfs2jn+3ehyPsKyuhEby+MBpPfpKz/5c6sobUv/1tJbCOpuJ4k7qmyfbPpOCD
behbI5guIzErLGhoTRClcH+CjPN1gIldfhnzy8kqj5yqmvaACQRwK+lrHMgFHm/0Rr6zJajtSi5R
YcRTQ7MaNU1woZSmFOP+wPQbq7HZSgUCaRhkNDCVu8FxlGC/fGksQiVMFGydzArGAZMLyFNMTJWP
Gq3IeQKqZpix4NlxRROjBzxjiCpQfGuTZtzMObJwgt6rqEFplEVBlWTfdFdK9rwpNGAGG8FffD8e
j4zAaxaYVWSut0VLy7aLTBypC0Pwsq/mUZ/dbcSj+sm66w54sjTypM3rK8SIMFAABBrBTOahhJyv
vqpWbfIqBNzBmhf1JpgQhg6s7Z4qdRMkDwaVtpxWZbMZqRuZG/VaqcDndSti0BeSIkYXk/w7Y/+W
xJc3vPALM2gqXNBG/8u4Gl7zZUAX9oM8bG0Xi2cxbgvInlsrcrAtLx9gRdnTziKKNN8B22gOM6MG
1N/1cVJMyqsnXTFwoYLENCxu14C7d5AlanfKzfnjk6/U5+gDbRyudIC0Zp88+/uTlj9rR8RmRz+1
40BFFmYustH1ZHPDzRxUN0p9nX0npLyYz/4UUmB/AmG3KZVFCCCPzANbQLbYIMqGIm2E5Z7XLmnF
iiXplQcgmTRivoYtLEDyOhuxFGhcxE1LELv7S8tjuPuPptSnyxJOXuc30DacmA220Ns4c+FReRbN
gdNAuIAZivia01Kcy0JjsAGlLqrTpe+B8yJ+d8ZBwl6pd2hcDriDieoK7ji9KBERRt7dZJBQqFsq
Y1OyxUeGWL+cCslx5xGQnkSs3aJVsttrPIycNztB4/zLZMattHeYFi4F/OY868o8k+9N/nIG+dye
p6ujmNdVkB3uM5nGIeZ0PKL1XE5T9QFM1MLCZkV2T714t/XzU72QpQZpx9+8v/Ex4P8ZY5gEcl9e
e899Ry2yVO2x9h/LSmqFyioZc6XeSwDqSsYJDniBZH8Hgi93wn60po0dyvHi2zB35yMPGJ0zetdj
yUUAEg28kG4DWSf0RRyS76Emd3wBruzur7JxoF9o+Q2LRC4F0XQ32KSo/1PbSjSOhLBudRZyNVtp
DDLunD6vAHkyjTRe5+84ySYN+MlXAwn2w8hZXYITE5VGnE+ZGf7nmo+yjyd8Cg+8Q8PCyIYBUG2x
bf1fdWL5R7pBj3zw3on7Dka1Q6hDvs5yGMfi12Dan2GDQAgYqWSKoA8Pj4AM2o4BTmg0c89zMq1a
DDCFBdgJnwazXprWL2Nu/TfFMj3f0RXZ2uE4YwlNsf/D94hcH50C7ByqV/L3ylZQ6GQmmh5eo/jr
TKujqG6lfmRspOU6rvKdKZUuJx0xwzV0mIM7yi5hlQ4KbzQucAkt0qhK04l0fTLOj+CSRWmpirB3
lZPaUnL9Iv8Y4vtIgEpN6kddF6dRNUXj2HW7Orabgn6GmOwBgsYCLtMUaw7bMEEcddUus/KAh8Ie
FsNegmgaNX18vTqa6l9U8H6a4IzPo0Z+AP5XwQd6Ddca7YX2I8bkWMEuqx/1oaCrfZFdDtJgdO4u
lkstzsjWPKTPnrS0XiNuYSOW7sWjUSgVdg0xi1zS5wrfdQBywyieyNAHTGMzY2qQuXt5hT2fSeBv
Q/PneNpByVWYUkxXUKwn/+bFj4RmJd5hfJauBkr/z4Z5240TKK0br3CMsgXFq16tHjVZx7blnvXZ
qrJdo0Nv3JG/gGGjnzdqCrc/7W+M7Wl30fWLQpq5pqu90znJ6DGtyeawVvPdEBdTDh7hpdjoN+31
PXEYCLgxbIlS8by8UB6bVcj9eDhgBkHM+VvGRnXwWVNP5AAJ2fCQGPXwPithdqZWNDMWsgw/RXJV
a0QXml6MmkDeaS+0SHvJM9y9BfnzSByQkNAO+PyHbZX20+rUMDCFWjTTkYQrwYbS7p7XUowWk5Bo
1HtjQ4rXQ6T7D4mwOFtgrzCOXHLRzfTQ+5NaKtPlGfO/BqXGnptECDoyIEDA5jAp9hOWaDjHXlYn
fXICdnNmPBVxtE+ojn4B6wPGXN4r5t/BPo9tG4SsmtuwAxUrfVZAmF6EcfG4Atd7vSNjylVk2jlL
LzG7bwvRTW9PK4jzytaDsk/3QX1Rfe9yQqLFVY/Z/dLf0PJY99jf2fKTRkSzupmcRO5V5OYr2x/j
wCIeFpyM9T+KbkCGCWYtBhZIFM/WXh5sSIMYZNYhs4x+78SEjsB+qECf34Fsy3akgkTEgaC9nhwr
mgCkPQdqeP5zni3u6tKfg7y9TuyWvL0+K0RJ7rDlfPYUG9+27AxvZ3rf7+s8QxkFw5rOL6I78l+v
l5SJyK5YJXEtLE5ldfnPJRKmIsLZLS1ucspiVrdZw3gC/rw4PDAYgk8SA6e/UlJsM8HLg9RGyN+L
utpL9kWDXEVBp/65NN1WbM9idAofhyO0L199JBiLo2WDF4bJNVnh12Ig3k6JaNvNIh8qqRW89IcS
qh6nZH+UXGSumCg4IFBaP3u0s00ysfz1f6V6iYAMkEP96GE0riWQwZDAjJTl9sDrxneS60AczbUO
lRIfseG11sROpAPFVfswBaoc58vJGWuLhSgk1ZF3Ev5K81qC5N6+T9LFhN7rBzUVRktIdwr0kBng
OH2y6jJp2VAofnjUlxjE9ooT+tW3n/6qOhY3hMFqmy55mUY7BZF6bLRV2FIGaCwhLc7M4bzMWqUI
P5acHtDgkCyrvAWtxdSXqjzqaOyDVPFsXZ6KSV21h9ppuNlHBnl72lJQaxvnZagqUVtaRUz9Z2FK
+L7OdwsPDEDKSMjEEPN2smrNM7rI9DMCwlDx1wtkncR0QIDZD+aZ4r2CoQsB459Imda7mZc5UMf/
yAm6MsS4T/RGv65C+Ywxm44FN7pLhNFaK4O+9H34HbTmOJluRzp2vmv9ArcEfynHTGqx/YhpM9gQ
t1hFs2+QU5hsSfXW89DBA4YNnq+8HRM8XVJ6qmHsKnkwz8V5CeLcP3Ryk/nnTvupkrNs32r/y0/n
nSBCk/jVxrWrkV8x2hymUXhhLlI1dIHb0qKIffn4ZYijPNp2h/8Oq47Mmw5b5ysGUPbjqYbBMexJ
uFEJdAHrfYo8xtTu3Jo8N/tF1BTd5eJg5E22raLkAvEp+MlpaRQ3Ymf0aYcHI7Nm+ZKeU9exsVxP
VrtrKkwj2E4caTO6JNHvK3hBt5H0Zk9865jcc+4CuyCaDRzcD4Hz6TEzkaryV/dz+fmA+qmMvCcK
ONnV3f+D+Pq9RxnVGH5iJlTwsvHlMofiYTtnyubRSP3JmVJZgIRqR/3nH4LtgKN6Pkz556cw83B3
4ydtaJ9Wnfqoxk97q37D1OBgLc1qyRJsTT7uM2Gbn+ymew1ZiIdF3Br2uZv1taWkdoLOejcGzyJH
D7cNuVnsUH2Q4fTP8gUzp6LbxQPihh6bGaTD2aJz7trgW6YJ/6XCIYNeDNEM0D58B9EWHf+C2r1a
AExzomGGpAr1hWI84NORUcTh7DWgkfrfISujDC6lPDBgiSneNyxrB7wDhf4PgbBK09hxJK66ISe2
Fp29zWSuRpuOTAEr011QU7IvF+YykV5EJ0AAvQGHXibjoXLVGlJVTIEBZZ+CfHK9tZdfT4cPQubP
JHL4Ah2d3hWa9m4dqaXzGA2IpdCLHYBa80U+PpYCLVCRK0EyExmo7dlllRFi1iAbj9XTltTDp2RZ
r7PjV3WTleacZ82hd/Q4HGP4f/RcXVnBF80BPkEZm0cjEAxdU5MRQoVAQTeBWXzrQFXVtJZIHYpW
IBtOTGOIpGbV3DsBLFvd3ki0WQ4GPxIkDAS12UY/BGWwwiUIWFtn8lFqCmNAdKTm0JfajHHc+53t
xhWyltSjipe3eFkmtcsBM7j0qJi8axOC+cY43Me48XhFTRyaLvdI2ltZpV5GSw7N3caNIBRADP4/
s10SFdDdZg5il7i//K71zh7vTJpVZxF5Ndo/zX9K7RVgMLj1pjXfTShNQ0CF6hzQFae7lXj7BW6s
7rHSHlGj0fvIXJboRSvtX4ssmbJ0iyd7A7Ucn/GCjhmn+JI/FPUHHhxCWOyJZ/mS2QeQy5mexE8U
Dx1PDSpMzHungZe6tpDtCzwUBxWGF0X2/R8W0gejJulAqKGgVM87zCSRuQmWxj+qd+OENjbW9au6
EDbdoJx9wh33MdBt+EddbgvygVQEf/vzgWx3ZB8miB0TSXs3nHuRiFAy5GwCNOflzodGK3hac2tw
7rsPykhJd52X2EImoKBsHKfxRofx/LAIS/Sr0tZDHNjjm2LwyOOmC1seVbaBloQND8j+kNtP3Ubf
PCcbaafxeF6IpSbDT2duPs7py9EkVdwJb4Z3nnznooiQuqffkcQX9dl8+Ht+HZPTZiQzDSYP4NWB
aKOc2QjbIuehRBjYQBe9x96K+zxICSbKX0iFWH2DLcFrmbFrI59TOSYHordc+2GWahK7dGFtOstC
fYOL7hZSisJsBCtZmbiQLKwTFrt2u4PkmLX5nBEY13aHlk+hRxETf26eN8imcTG/5vz6fERO8XpS
8x3OIWpbc6miwrpWK6MHZI+b6xLyj4RG3MXrqqzpLUKEPr4YDVl8gBLK+26GjxS36qPv9kOGP0LL
vfb1iFpK7MMCdZj3SlUXhmYSt+1Sa+vP+bhXsBFuUDAd1MhAK+GdqoL3rNsDsNN672NLVfZ0VctM
mmJQDrFXQaovYNSVS6bQcVs4D7OUdfFBRO/aad+rudMj7uoMXCEH9cVcSrU7W8K8XpcE/C3kF2ci
wInEz4kqNGAWb/dpAwfySdC33nS6L0oNF0RqpdAhtdGJayjA57230TP2VTNQPMpnRvSEBnbEo4vf
5O7Tz1uTQlX2LKSe5p1PRgYBhQUdc4XhtCFz1SYUH1qXRbPPEo1G+BqGV+zySIKrJ03tZRB9yZnf
4fpK/1NP1d4T7dIqnxoqJMw2iMyLt7bdbrT95Pn43SI2eZRt4R66dk/ImCxZKNafBYDGHWWDRIy8
DmR1V51Jn2GwfE6fFFADc6QjgJPzd/66CN9Ahkl7oS50MnmGJxG11aMHwCUfGwYqLb4heqTAhMJg
4Ragw+RaHXrF+14uvqG4U470Ax28/9K+XaZd2M74Qbj2N92PYC++NNWN3Z5WCcguFTmUYmzTsfdc
hx6AqcVWe8xsT+HwpQhapD6AmtMDjcKkXVZNKq4Dn3aC4xGDzZPxDwCWgH0fFzDgHdK2mSf1FiQy
GcT90WSTi9CDvEOEvKdI5QiyzWljVGRlJuteOtXb7RA6g5gyDCZ8aAbkY98H7wB3yf8Rmaa3nVak
OiR0jpnWioKwTJWHa2RTum0TnEiMjFrTvdjNJnEO89PLBb6d/JyNG/ap0AKNiBiQIo6GYbk0HJIu
UZBH224LGiOTYzxd7EV9W2cI+xD5zQxo4dKYtLPZ6VLTw/04wSfKCL0C1igm2QeWDvR1Chxlw63D
nF7hOVUFyibUbk/JKoZCjf/zW9utXt4P7H6mhDGmo18TiOsnzWTYXJuFA5UARaGVOw17Qt5hY75l
1qaWlGegTpoz7yL4NSHt50vV5OPi1YGBbZ/GmnygNuOKUL8HnkiHSEo8Jn0lerrC0Dg90YxxwdHY
IIcaXQcOuxIsriKhfAXpSpFFs4wGIcaNFFcexj1BgJrW9P0qYbkGn0SuiCN+SxPB1AIS9y7p/GZf
XdIyrnA+TrM9kSUyc2bbGVf0po44Tjo4RUu9yg1W/WACEhnKaw+/GdroDkYN8tSM2VE+/7I8x4Vo
mOqBFQpTg1pT1u6dp4hlLZ/ooMXhoj1Jb0nzfjLuxTSlb86ORAfGYxbbGdKDvJwARQdg7i+xaW8h
GMxpRZBm/CpaIFz8iOx3nSz8EeLkD9g5GqzsjvUihpJghNpq/QlTcoxJE7gtUJAKyiDyEeW8DZdv
CgsF48TVCuRrt9fa9ombRMTjfw18K1totUvFUb4aZx1ns1VcvoqHf6BXeZZuFEa1OF5HKFih0p3I
bC/1i22j9+SadbKgdxYkRQTVdinD+IzZn7IZQSfZ3mUxElHNqq3pGrSShwwiySqkMCjmms+HxwGS
lAEOX7q4Aew83jzNPm2PfL/7CyVYucB/7JThQ5Pi9EQp/WIWGWw+jV00HcKwC5qFo9ioOkQvqCrO
fN1CnUd0wirRlWXMYyr/fxPRiSA6Zy8pp8OT4gwPkP4WaAVb6wUJaOVANvzmAcsoiucEma7byWCh
Q8oQEAVPe0CMlxjbCCukk4dilyZGfzonxzQuxkz19IPBHct7+D6Cnz/ceV+20vqKqHOydDvHDGoo
suXYyqIm8bda9+6hcUAJUATqOBothW7J9EfwREs0cGM3VXX5JXJYJX0i2OWVyZw0P4ftPZS4jyim
yfi73cSJtwzN4vPe6UM0zf+nZ96hGDPedjs996a6hkz2QHXe2R4K2y62Ax4BFqp4yCKumYoHisDX
rWChtZOZAM0kjqJ2tRFtclKu4IExybXu1E80T8FhdKe3PPWd9ySafxILRXOsVB30XADmYbEPfMzW
tIT29YM9P1VhRi7ayNxkAogROue7hfXGm3gR11T0+h7JJabYb6umRM3duPyqB+rvW4rQq/d9+PBY
SVWYF8Kog7Wxsd0zeUxbzN3IplkxeesCW1ZCb2UeuBrTkpUx4hkmn4mrRfa4jFgg4Dx3TcNpTcln
O+otkFOGi6UL4da2yY1BvO9OLkK15V5DdMVFa2AV1xrMhbj+k6qAD7UnBAUSEk19myqXorKADEQN
1aJgUD4moRKO1kHW1a+kKAr7cDGZenzuwxb2Su3enmicnUS3KD1B2JkbD2MlP9AXLkmN0NCYKO7X
+nrna9RsQFHsxzjPZ7RzRH1V7/HL/CC9i+wdAUhUqw/9tc+QwB8zwjPF122l3QlXrgfInFZyTUYj
X+7DVw7A9DcFFRAdoFvyrIv1TXmTyEqlbKJM2iHZhWkhjShJG7TzERODKKMQklboqNdQpy4IPXr5
DHqoiV8HV75lGoWkfFSsABzQ+d93GAGPTd46sHs4E2D7h/y3Tvx+Soub+L2BqIhIRjgwKfOMY1ph
dlIyH0yrhudZ/pbG9/E7tLg8EQi6hKFOwM8myktFcfKyfM1IdbOIOaiBMGmd+w/yQgeCcSHcbK18
H59bITLfatDMVUFVbRkFy1REAY9C9OgyZtd5L5amUczruhDE4o+XwlbTeXFoBCn8YBBjV3l5FNJu
Cujy2KU2jsYPd8qHipuEOtl4S6L3s5Fgb/spLTM1+9SjyTrK9oK/J9tchx7Nk86tCrvTKpwk2fdh
gkVlHB8wvcM/p1Ki5b6brj1NqdN8/CEbY29vsJJrlRjZhp0sroN2t2DSD337SQWbBX/q0EiiuoKt
FbrPSjCWDA6QUQIeu4/NLpjuF9XOmJKMSNcuGLRruU3GLmmIqNmofbDa4HasJxMBT+lNGNHo/9CD
lw/GHQYSSEWl1NYZSz4OmfbzTk7Sxy9sWO2kzIWcwtYjSfbk/O+frVLX5A/25797nBpw2Y7+hbuq
+XHge3pIjfoknEJsEaDgGBzbjNkz3XE0uC5bavOfv9m1tXi3liw4wjX8teWf2PJD/bl8qHfJF5GJ
U9EyY6h7mSMQs8mAbcCXcIGtQ76lvHGQEdjg3iUpD8t98zB0cBldxWLeltSktxoQ10vYQcA5/a32
DZYXULF9Zi0RLgg/5PjpjijJiZRDsJ5yrEhVtCJV4bs05UwH79sTQZ2EfB9LKN3QiAm2V3dhX5m2
xu4/2kMkDDOIl89z/wjKAH6OQLS4mOzpIfkaCDAOuBG1TR2IPO/i3iq0E7ec793Xkrn/Nf3ltQSf
ZxB2LAs7wPNzkYZdXmnzRqXO3D0aWMblpLdD50Y8umHfyKL0ZGNHxedSZUB0iUTxiaxTjXDsm0r4
ausdR+h9bsHcIU6ROJis3iKDjCG0fX9vg6P1C+pf+BZIa3xTdgNYCOar7/WMdMpNsOl0Cc2Y1bZc
103qVtgUtNUOjU887jsD1CX33ZY4vxJGyLgHw1SEQIfQYl7s4W2QNKLfkRVMM90HWUO+KpwEnel6
0OXKDK30ylodNDc4R4WCHGJ2DNlMEe9WDJ17GA3UotG3eZJ5eWGMAW06cMbP9+J6ROIfJTvRzcfx
CblPikYaWMHA1Oi6K5Uu6U0HjmcRi1xprhTTLECOSfwlby6kMVe5Qib8wGE5YyXmVugqknbcLFdm
vcHecEKxB6wEaEDoZ7m90PmN/iGx4NgKUvWgQc0ovaGTfeSfIy19N9Uy7zWwAMxm7x3bmQKK78t2
bvA5rFeiMCafEnAA7XaJh8kgwL/6lzHwPF3HrHmFS0iqnu+kPhnf1ms8rR1ieT45lIsip1MWmsGW
HZ+hEjqgQ5Tf4e0XiNfxOAURQqKCwVA0mCntNPUeHQTwh8VgafeeOnv538FEHNp6b0n4WLCXa1wK
/2agSuIDwmcWWq4ZMexoD/3EcrG8VybpKwcShUcxjhLBYtPIi51dW8tUndtSg/skqAg/UjF6fnum
2+gBjm3nOHgcr8mVSxzUirONVvJKAhLyc/Y8OPX8EKfmHCDEFgSGS6GUAQLweiYo4BaQ+ZS1ydlZ
e9QWJI1QJXd/p7b46cuXNiONhlPs/lr+PITw7BGgYzm2TnAmkASFrcg18CtGFm7Y/Xa4H4RxtWJM
BF26QJyQNxDbgUNPseNPd9vj/RES4NO58uDiUyH4oGTHhr82fpaEJ7+/KW44d34TSfXwDLiGgrX2
WdMUYyXtRgKJmCwfniq3u5i9LLWDKhkfZNgi8bbDgZhfsD9BGLx6ybKWwpj8tRd7H7o+i6HOYwcN
H/qo9ee00EPMGi3Sk92bowBTi24ocM1/fHnBkduE8KppRVS64LcOkAvprgYSuwEeDBnrDs4xKA6A
+wAOo8t5VUPFRi/lKTgNwxoSAKYip/bU7hdH3wpYnhuX47X74DQPxrQUfKhuDGtYB5Uib/4STzN5
9GF4q8pBb3lI5AJe1egkSxfRj43FDHCt0u7xwbCWijZoblKkmBpQCflo25NeeR/kVFaBvloYCuW5
pRcDMtbF6QgUhx7buVeuAIeV1PVGh4skv/T/eQtX2+d4s4nfkGZDCTAt5AJbcv/Dy3NF+QuvJCTN
NPawF2ZwgszmZAWzEw0yd+l3WWTxV7Kjm28pl+6DzfBZGWrJN+NqcZHrtpn4jycpxr8GYp4UbHJv
ziU2VLbdi1vyp/4EEAAZn4zaDKhPFPgc67IG0SEfUkR2vTVsmsh0m5WWGviJ9ak+/Itj5myqUuiM
CRfdFVCk1tTmBGe8CgU9yEkJYBiP9bXdZKNuDPyAWhGoK3GQeZw3w/6V7s/Hums3epv6fFWfYrun
BpI51CGouRS+XrcVHDUPX0Wr4JdE4Q56nZ6R1TH7Q+8ReqqPYFJovpwNDLvb6cPY9BdQiJuDsuqR
d3an31jIzuWdluWKSQkdkK/IG8x0TRdTZeokiru0ckRWhEj1pTZRfHfQjk/2p/HT11jymXiPDBzm
ogf5SI8EXUFX6mGeUll1P3ccW0ZHbT24NQl7/KNO7lXqPyFB3TW6dTPbeEvSZQ5/2EBej8oVy025
/OZCA/uf40KqHDGtSlHePK7B+vs7vH3yLihwZlzxh9cdUgpxOBMy3cCoWwDu7CRAdmo4U6aEZiJW
GoW6tpqLeDqZrk9I5WDlOdW5lpj3dFkLjC/O53DF2D6XWayQY8ZRKQnBK1vG7if96O8X22BSUq8T
oq3qR/2//4cnyb6671HK6i7jxOSZ0CI+DYfWl1BuIj992TTn1iaRzYXRgdm8lkHd7qcw/m0hUuPh
xFDkAYQpuSvyPXy23pgB7Ck8Sqsz9gcvDseBAEqiRFyRZDXhSyanC0aeImUSqrn33QPNVfZ2oewo
WTv9tazcG952DfXq3cXJ4T/2ipahArKebo0W1Lq69EZTdiHkV8zKpOIYu0hJrXJmOgscNy0n3ONw
8ZaWciCWDzg5iYbl7Pgn1ZKkKVYBMhHa2RWmRs1I3zvprfuRpMLy1q+z/V0eNwUhsqzmdpnLCx9S
KNVUczpR8jS+a1Y0A+hjoN6OUDq7ka8IthsdKYsTizzlxVShc7YZj/k8pKwN8YC790b1VgS8zmOQ
o2kCCECIH8Bc6ZmRxSmnpV3HaplGudGO6A3rffWGfkpi406nsLTdEa5tPTIYT6sAHzV43Y82hGxa
TlVpNoLx/9ndWSVBRBKxZMyUQVpJR4+yj6RJ3zHlIwJWPtH1YvFVxrdv7obA8a6CG0fW6sJBO3+a
FaJyDPlNbOyL1ZU3o9DZgefk6Sx50DSdxEDA2fsA700oaUQbbgV95TyDcMfYfIQCVpyj8biTbqIw
MWJ118s902GvQS1+/rSwpy32tBvArCUvA1tG3F+WEyFODgMEapqp9HEX80Klem0Au781Q3aEqTl2
9w2YEHYcy8Frlfj+xniKQjixYt7JV68OxveHm9QRPwsoQcLHjjQobFgAWLwG429ob555iDbunlYB
x5/JJ+FPK70jld9J9bvGTfNgEl0tL1WklC/juqFdly9urFf8pOG0O7qdyDsJhBEm8br6kwe6tYcm
/C+DKq4jdPIvJaLaPYzGv2LHXo7lrNLzazIwnC9R3vwk6DeZcKMhYWIC/PSRsA2TySjJKoui69S9
nvUUZ3qL+uqyUk1lUlEp9jKplsQa6IB+tAdnwOSbbHxW6HYLKi4G9yLD85lr1h2yRwSxpa2VsFBx
U1v8+CxnPBv77TjAibh4UXnafg3JNWL+XP4NFLU+kVCGoxMYM5nqB2dAviFVzb+gzW8FVYDgvCen
g6v8z2HFYHtvih0BIaCR0ZuJH1KtXiPQaRBgW0HCaOm8XJBHsxZcYPZu4zT0q/mJU/v36WlrPlGJ
VSlvEDhzpq4rEkOuwHp6NW65zp8KTc2HtC7FrEYu9+RRs8CQ5EF13hMVTdFg8fYGgxAcqgBqGEeH
GM79yuRQl+B8SU18+psGDJnmsvL9opeKZd2x8ZqS2wwmt9Id47wsauyEgdWVvVJkII+7+rLoVlAD
px4WB1rAXg4vjgYxW0ozTNq6+5KzqCxSSDKpiQUR5NrNiMk/7Ty1kStzHcVRdjoiVnSETNvIw6fK
PA82NNjkPVMo6sQ1zSuyYnFx+bR8Bxr6OZVIxewlOh8xcZz8qq+G9s/wfM5NlzBZkzQVabV7DDWE
0QbThlQyQf9j4Mp41KCv/9FC6x88dSk7S3iiPfG3GBEOhnuiy2IaipdK/GGLwc6xhM2fyGBAhILi
kwENx+ftJ+tCydpS7Qm2Aup9hzr2y5BSpJHiQU2AxRZwQ+d1HWFVGO7cf5hLErujb9zBUcm7dWmB
txUcgtMmQAdzDN5Hxpil65rpQYpHB4xEvtBzaIn4XNvPeJm5WtskHN/Ao/5teWhLozQnAVXG/L+S
s7htlkJgXqY6QAnXpSyVv3Noagq2SqBLWk6a7uxGXZMNsCW904R3LU9UBM+LdzyBmAfNmtRHBCrz
m40zvNXAVWjWe+8BpqoR8kkVPIDRuEFJ6Axyoq2+ELvs/W/elR83wZaCiPmARfKoDHM1ZGn7c20T
YHRzEq4cF1I8FsCNcuq7NDNZVVwtHd8yqbFtKNt+twtXV1NsFZmenTHB4dOEI0+WkbMA2xIshQhe
az+gNOic1MyVy1JHTS5AqVWvdWHe96e0H9AwiI19Y5tCKYHWFmVgngEo7MJqtPRSikAGFJkJriFZ
fQeoPM7L4xRPjtbd88RWznuUhtHPOCQqA+KC2onubehFJUV+YkekOkInxJH6J3tElV0FroN+m4Qi
xTkbTl1/L7L7JJ1bUaQBAvI/ZbIj9Jfz6otjfgY9NOt0uuB5zaXN9V29XsveVD8TIc4NkC6rTuWb
o9X1jVZ9KpyUtO3nTNJTis7ZpJSXcYMCn+loBXflmUy78+zWi0g5nzJHuxTWtyKlrfLHSO5JOfhB
RYa4DY0XYvb6+bYp0qCZb7lv+G1o6NBi5wpRFVeYDQm3LE14jhXIlkzsoZuWS/hC9RKWZLVDsQh+
rz7tP1fZTh6h8DTOK10kSCGIvixEwW1pE0OoZs4YShVZUqGs8XaYRamY7JgndKJpJ2RWvGexpFrH
HWPRhp/VwslCnpnNApO1zuEqzajdzlUKpHw7eGp/ZIsVOZ50tlf+RBSy0GaluLMdsJIufHUknYpj
iC8ihNMHLsZX1JP2okI347ng4eNuOngC5ZcjzMOLN5NybIjxN8iZL33vm7tYjePuNp66ZVfSPr5F
oowfxtBbqOQH+AaeZtPN9Zr844RqqgZCvPfvu+0D1csuC8JLySabdeOENlA/v9xJNWXac4nyeT9W
Vxjcp9ZLmBq484aXjbidMnBbFZ3i88d9c6PqrlicawwIjKONjDc3BoBjwyNcqSQcKPFnPW9UaYtv
LCa0K88Q/JHTBNqjUmSkJpNssBF5wXrvG1eAnKX598FVkRfZRG3gBry5A1BeRs0JYiFXuWpxbajv
emQwWAelqxQNN+dMsbZ9VwGF1O7EW+KTz2mtflipkQh6z4VKYbRCWgmsCRxiOk2mQa01q/qW5K3O
623Z7eFfzm92ocq4y/SO4EKUQ0vJBheNy1IpjoER4e9kIWR7TGOVhkcbqw/Deq8k3N0B9LbkK78K
QTEQ2kxeiw7HHJQdL3A+w/TXa1h7cOCYXRjXCjok4GEfHsc+ctuG/umGA2mLvXCvkryIvD7J1EB9
KdSwqo44u6xRAy2K1nl4g06YLhCUefqHUxIAcR9L1MhjsI3o19wUQcu5sd1NTJ+j9kRFrvGoK8K4
GNUgdtg5cS89UukfvF0HLZEmmOFBTaI5ga6/tWN3aeOeAKN3jVMaFm1rC9upESRgX+p4sDXRzCyy
G+6Xd/t3nzEjityd1goR0Sb6OWEVJX+czGnV6WT/XnvpTP1wz18zHmAiJ5bp47mRG2rwZrpab3he
72NZws0eh1xlazstdQYKOoCWE5lUtljdbIxjssrtWjz0nr+/HHrNaCMSELcDnMrkw404I285wZEO
DQe4srDmxIQXx5sYV5HWR4ztoF9w5H6x4D3S4r6XWWFSS5QRm8OGawdFghRxvgWDJusbMDsMzBHB
ZihMZYsGQNoGUR2ecgzgJG0m22iuEOZtNZ/PodvoTJ3ocihp3LQAEskyxSqHF7jfEWdaNYkHhtqu
GquojzhADyZKkDdFEvYBNfDjpp2nvquVbSQSrLpTD9hrSu/HX4Wz/U+JZNu0IppcDvCV8imdONIh
1rupsMq66QrmrpauYJqr3Gl+C5/SjqSewydXJJyPt4rI8KF6bz6lJDaNeTghXjBOAwQEMvgkl438
1zR5kwAQoZvyGVMzFw4QhjVouhlEU2J/0Szub3hML+fvTsMfR+gjSjGoUChEMuFZFgTphdE0R8Nr
E3ezJ/HjEM3kz7UVaC90bFDFxeznpqa9aZIej72bAAZgm/PViUbr59L6gfSktYPu4v03ukfAqPUJ
ePSfnFe3/dIdSt0YMdZcJujsFeOASA7LOdQJm8y1kNHkJEFUttiv1tTTVXmDDY/A4RnSDhcMz63N
v7af7q2dJj3579/6xhxuwtOM6q80ERyNP1n6CYXiFkO3gILK+NlsqRGry9KLWAWrUjC8cAktr2m6
wN+pFtG0SnpDxrfrJ9ARj8kw4QyBxx+ruTBl5e9PvrXsjSeSUB6JzB/j1Sh4abF5ssn+iWnGM1jO
OjCfcTJVIAOwP+jJa1wWOezLzsqFNxlAwEHxD52SNFPvNn8JS9S1vVIsqZ+Ck5iuGXHYRnko+T0e
OQLExpqG51GkTQWyYBQdTATJ6T21mqs1fzejAM6EndBryEQ9weuTuAbU8PUoIDQpN63QCsMIKvSL
ilvLxlNJbnQ6KgqJKCkvP9/ykzppc6GDRjArno82tYA+3ZMJ8yZlcq3imbbTwoK1ZMlVz3JqjsRZ
eMmcwrs//hEDOONih39+dngfGPNQn2ihwKJjNJIz63KJQqxQhSiaUcw23MCR65drZnI42ATZT0yb
Bn9C7VG+CjUp165zJ61DF++7kzDph4BDwVYjWbtjyn/CDA5kWf6oL992LwsvwhzkzH7WLuy5qMdW
endYkJNS0RDc6z+h4ZTKhM9Hwqa2Xt6BDLlaBKFq0jNz1nxpDSrAIWRFjUB73r1SsFhvLVA/0p+K
k9sU9xQUeXhbRHi40dVtCm6qlBG17mgDsBUrKJRylwjNVdyginfgCJos64t0j1fS683nyWHzdh4i
4P8ciz8Lulq8cja60Vqqoru5t16YNd/GZSpJnp0378WsdRAmuy2S3BF0BsoiBdbp6H9gyYpqZvUl
HvppHvnz2ULHmMX9rYvCQe8BuX+/jwfGaMiVQ0gBbV4DriiiFcbqvgu0CxdquAsu3HoFU6fPMHu/
PW5iuypoxP2ClijclMjfSF3B9HhtM4aHj2FoJ8T9pKxl4B2Kv4vdtn0M7cDk9DDcnCFztsEVdQ8X
ZLZQ9tK7UTyz/dzPTEoXEQ4p+dh9Wa3in9cNWUnPic7N8hox3sKmxbxZo6dnt7nWQHFPZgUtlNuG
P3W4ygMBhvsMw+m4CPKyg5B1Mp/Rk3KJ/KqVD9msO8VniloAAq9HcPDo6NYqF1DlwqSK/gSTkZ+L
oCHIttrRbOIiX7YyU1upBxm9dXQNDXNqEccGYcJdmh+O57zB98RE2vozlDYztJbQUGNPCp9F/ff1
rrqZ8GWSUpkODpbBXAuQb4r696tpis6dphXtdnuuGovhDxDPJH1D5t7na54ToMgGPXJYc+FiqRfR
oKFFQ+vzCWCEpDovX10GmaLDMuZAwUF8VjBsnhuZ7FPEWFcFAkkGCwz93IjKQFK35U0rsVfrq82i
M3Lb16U+aHD/nZp+z+govEDM7Hq7q7SWb5OHhI9NgKcbuLWma0Ac/iyrtPMJ8tfZRUJmf1OLrVGv
hR4lghHF6FRugMZjXOgGnXi7gMw1BT7Vq9iR+L0HxbnS9x8FPd0IUMdeKIUUzb5lHf5Obt0f6lve
1gUI2A8nzTJCP5viGQsBfffGFBr2zuCWhAhUcC/we34qwkt89h71NlOLe4botBOkrkdek0RQjiTZ
I9x5Cq8LtR2vevJIwpfTdmsvxrdAFNmpWcCcphKHOr+tEnIQyUAYzSvJsa8fa+c9A92OIm1qSINl
1IxFPkwg+2AOIXs4CFjPkKBK+794i0j/TChfVWeCiSqHqsFF32fwg6sPl/6C5jSbL2tQhUXCVPrb
gC9gIuvCfeqyXr3NXv6Eutl1J8o21DRMXxS7kzkH4NbnNTj9me6PHhUM7AubItjhow0k1Nq+50Wx
yWpJHS6COUh7f68FQjGddTR9sGvWNF5E0qBo/tNP8NeBO1nczv2INnxTJigIOF/cKed7RuzJAQ86
UuCZyQljMgVBNFGWylEn2TjMyksvcXdm6D3QV4FLW8shRjQ4Feu5T2fkT85ynBGW7hLw6MWsfxr+
irUHbNCu/tcZfOkrN1mIctrsx5/vdvx9yIqtT4Ypd9K7UsuAhFD3RzCrOMlzboeptSRaaUlVaoui
RoK8aUISLkVoCyr+bWIEqyDjMwgWQMQ2NSqkIjZ8NmpkYItyBDYN97Juc1zgclA4iOFeN7JWf61z
TE56wSi900tFBB5PA0n36/vo1A60xFURXpqwMNc5fkNld5gLQyy7cycwdqrJx5f7ermkumpsX0/1
oqU3VksSRTzMYtGoBET8CqDMa2/B6t/AlMdUt0CTrCNtyTIvvkfBUYlmutrg5e9OlCDEeBmlNiCR
+k3PhKWuo36ZkikU/j0TVskz0V+W04k2OG86jGb802CYr8pq3DIbcmMm3QMsXf4W4z3CFjlylPL2
KAsayFCQT3yY6fDmz4dHi53bEsWL+dPEJ2s09N4L8b6eJlsythThJHHK6dcXKkPYqmQ50weGd1sw
wnb0rpHcWfDRrtUpSyPPunfASsA2uktdrFqV/i2I0MWL1MxXmRz6J2a1fzwkJQG7Amj76f4uYaFj
K1ZLZ5JLO7BZO4rEpL796S3naHrRS5xEfFe4Z0sZq2ZKtiYos0RlXuadSn+ic/+ssXjYLnqzoKnv
mnyd1Znn5foLl1Qt/Q0Rlm+pgbb0ok11708okRYcaayUvQycCxos0RuCVP/fHyLNKkMTrEz5HN00
aNHlre+lK8G405N6bD4OClM+fMQUzDVyuogn3yaRQXuK0Fad3uzZAnp17wBzsUHBxoCo8/zXzXYX
fxWNqtc8A9AZad7bGQeELomWGqayjVmzEw0hFls7T9WUaa3p6QXwWgvIhHvrWQxMKbqNr2qcye2o
ufQp9pE3fbwCzvczrCG9FAytVXXlY6DAg550ScNWdd2QCMEK2U3os9lKlaLEpbvA6bww1EHsp5WD
4THD7SF+Hj1+LkbXsEp9s+ssTzLJoTFSSmi8uG4BRLWnNPrjQu9avZg/jhZfuQ4mufOcFOl7QZfU
InG0rJ5jjecVbw+0qy0w0V+/nkF7ZF/XHEFiuD8Hp97mJMjfC2IdQcPukiBdbQdwYzaaK4OTZs/P
Dt+FENxq2KnoV1SdrJZ8ad/9UHhtRV1NOl/uEnu0FQ+tkPJ2l66pv9Qw7TiQ0MX00F2KBfy1buBr
kxfn64yduQgP95zXP2ApRWdv3xlWeRQ94CGbqLbMl/M5bplNDty1nNg0F25LAwRkBkvc9xUun4EH
mqsIquNU5DV8SYF52VaA1Kdil/Shf3atpxwndjejRYTPt5lN+64RBND23IMPoUztNyu/nX9t/NdO
XTsT7hpCKm5foWNQMNA5JppasCzcFgBBxCzMOyaG/ROGmIsYL+NSsS/mCWBLn7Cx6//o9OfMOLwE
mk0oIleYLZAVfk4i6LNwUHkTOzrScBHfULasGChSfJI4yY+8dqdzxExfyULW4QSWRlky/KryTJrh
guD6Hzxk7YVpfUQtQskJwEe5XbwTSYc+12XqBQ83eZdb/Cx83aPykel1QUeyE7DZdXVQdw/gMmOa
csL7TIvDRw/v3gZYGEWGFNvtRK0PJBR/dpfmUMEOwiyb3rRSB/DSdjoH5ZBzdRyIJ94yBrax4yt9
T6wHaDG9M5YEN0QdJx2uye4hIGFRGjMfEanu1GC3UEwIX9rFG+M7xMhMXJ0i1amP9qGExUYAh9g1
/DtlxkkyiZTrgUKXWOUgK5FDmFUjIHyr25zCozLn2gj/bkh1CF9yYnNvbOf7NGLlVU8RqMCnnXz1
c+Jotmpne4qGLzZcWQLMl/7cARpiBYkKN9tNwt8Unp3qc9E7fvc85yd687NoOVqOjoBAJbAj1WwV
ky+YWCE1S5/RukgpJZ3fU4fsIwGJkpLw79L/uV2nEIiQT1e/ArZMxDEVHWLDJTSJ5czzeUVJ/7Uq
gxma8auP8PRyEaA33S0Mi7wwjaiSw/WW81YRvdCbAoNYHxiiqDsMVuXCi5aqWLReSf+pjTXg0N65
wxUvhwrUB8ouKeipK2bhA0aByMS0YfocQ/4Gf0bgSxLDuKWOoUurkOkonhV3syfWE6wDO/TxltgM
QI4aOZ04xMB0s+21Xd1Ee6PnRyvLvTGvvEsnQuzBxmhp/swcPSEPtXE3aZd5UV8HVn162SDEqKkv
TYIRewATHz1vG2+CZ7yPuP9aKW/JvLrkCIR6Xph4sWC7b4sYxyBcLytnooYhpL6Ypc0Ko2IgsCMF
9c+jCvT+wsUWQUxleQi7GQd7d3MUYOhaAunTH4ISAegm7UGxMy4DxgPzgEU+9lLsaS1Y59p4sJJW
vtZXvKFGBNGoZ8tHfRLyktF3ISiM0iMxJPag2LZKMWQcJT5dX3Xh7gM1s1goMyDiswoNjojFdAFN
8br+MZgqnddyPWVurloJhdyALbrAKlQUiYSpO+PUBmcMJZdUn8uJ507ulAyhBvLP51629eOJs3+7
dnVsyELFPYQIk64QmHFkayjO5mvHPOFbwxCDcLtwWIL3EBQIV0z1QZ6Q9GHGBUgf1qkIxSuFoQRL
gR3Gmr6mbWgxGNP4HHiApCNXGxD9Qh+UFMBGR4Sr7PwfEg0R0WCNpBmziyZtRWlz8A9UD7Lp4J8P
FksUcsAkyzGcQ1gTJlA4wfwjcxqX7qrgEDndRpzEjUF8AN26iLcdo/YTqWguS0oO0y5drM4EuzWW
QvKHuXWuyrx+6zJ5W6GYa9tesj1zarwUt8L6XMrVNsdrRV1lC2n53soEQmjAObIKZiBhqzsMUYcD
INhosyMC404iM91R2HQZau1+t1Ultf8d0F9lyWacyS08nMHM6m0X8wgdpqGLoFma6OnLaSV4JTuv
op47vs5/TzL1muYAUetJRMvs42okEiYAE1G2oArmyPBGPuUO8J0pEbJ7eFrPANY8LRepxpkUDO6g
uSUFNpU75y0ptpX4xz5FkBtFPV6NTHUxWZymIWYbRk68fll0nkVadyIyydsOt1FScBshGegSNN+0
jNLMsCtG+hRQdYcQj+GTOJAvEWt7L5tK+wWu3KBsuPnyUxDamujzQX4JKnjbL4agC7NNLFAjoXt5
q/yWDbmKJZQeSZhWdkuxPojd+8yaph1imY+cKIvOcnY4TA/of+syvG1Yo+gqf8PRbNdrV8UmRSXZ
nT7Ecg5CLp9gS7GrPT0G/AQB1dPYubCF6UBUm4RsQ7+zzyjhWtAItIUtcmt6HVTZAenIOar3uyS2
mxiX9LcgtuXcT9y/HbZbpdhr9wcqSIakcP6MVg99FK4Tn5Ap4UdlA4PRmyYUkax/GH8S0CV81pbI
MomYr6eqD4bek72c13J47w7m1zl3iF4G0P3kUcT+xft06hNZSTbf+neefBCWiBrQDF5sEFQzA7tL
nEIe8Boygci+NPcxwVFlTDd42rfhKcijiqH9jndW5mgDSV8g1BMDY8kHk8wJ+nEDTHIWKTchECOV
/rB6RoQz12dsJrqfpNEzmtD+WCRZkp3Wilcpd5mqkmJClV3eBKns07Ti3l9lQtsna9c6jpnH2sDg
vO95F5ixcdScsQZKMzGENa+LMwzlYbTxAQVUJcR+IQ4CP3XXSzKCqMdnkfCA3VT3C/arC7pT4ZZn
rxqSFuSs/MxtZvjXw6Dv1uuCmbq6kQOP8q9Msu3Uh4t0MJtCDVT/FBgk3VN7KX8l7BgdUfMnVxe+
g/VB28lqmtB+zwVyx3e4g5rgncoE/leED7SWlB8Szd0QLw/hVy/Db9J7dUTY9uzLklrDgDQY36g5
cnOTpL7mohZug3lal2AYqouorDH8gsdNDydBXIEHVB0iAOZEpcPqNjUQLJ7qUnk9zesyUC3TOOWS
ycl/cqX1Vrzjwaf8cUsRf/r13I3TEF4bmbfmBURFvhW6aKyHmkDh7dgodqikQL2Urja99fA6ddIX
rhtdJ6L6MQf8ezyO/arcRKiAHZ4LB2MyXTWgZHc5s9A+KV8bmIy3u4EIdkhwY+hrDf7ww/tDrKKC
HQwvkACcvFkgSzprbcrirItBszfyO8OgkGh2TRgrPLGcVqGjBcS7jVy5cpGZgN/9nlyg6LbcXDpO
ndhC9kXHTumpnHZuWRdCbWp9Hm919TWqnzvUH+xVcPQ3SFnNXtueJ30FFZ9sqMiHW34zmiNeVf9g
BPFSd2a9/i3e/mCtfGQw4bhXTwpdKvbSiePJ2vgzoiHt0PM8DA2Zu5ocVz4I2AH3PqjaUQJnPVRD
rUn/RmLZB8eKZQ2zkj8rkRydSyCkHvr7fgQMeOTCt37ZyXfUb3RlJVCeqiNEJngxp5tBOeHr1VfB
GOejSCS6vRq0NYql/3OmBbUuLaihNJ/LEODRTxcCzAf24Ysj6ubrnWO5jLpX5vNci7wa1TZFvqf2
REgzBQjX+w3B8Rl/1UEaDZXTuUSEsiDsqo2rB8NfZFSg5UqcXB20avrlWf1yDYzUr1Cne50XnH6A
rPTZEhcUVefTFJvmEPxU3cwNb48wzgGXCY8BrcmCwFNN8MF5KqtpltoLoolQO7fdWPn4nKhHqKFo
Z7qUObx6lxhAJoWY0Dl6ndqgxp6sWbL8AwLW6hqBVAjWcPpbmP7fvI+qp/o8x8e5YPJjNx/3kY9B
PGaBZhhbkWw1jDZbMBV6DfNJh8ay+Hw0KHSXXuXcj3TMoJ+F5zWBouqvYPB39CqXJ6OPF/CBrgXb
fl87nv+iXMFiDgCnfj7CrIkH8kBhYI1BSgQUkRu6C2S0Jwp1TDmb/MgdhLsb5ovMC1AW/7oYUk02
eHUXk93F3K51nhlfO1dPwx0G1dLiCxmtmehzhX/vV3pxhFgYz/E9ErZPXuDpbU5BUP9rqHUJC75j
xiW0a5ZV6DXB7b3GCpZDxFIKsnbj/f0VpP4hAtG0yicz7KQpHxCHvG0DkP5jvHfaw1hR/qvCUEJ3
fmWWtMEOa6yUYBWYCimQWY7wUxaSf1A/Kf2d1NvCIkNP/I9AOVysvEyPxR4Vj6uf2IaZUpe3slkJ
8kWI+s1ayxbKUw4076N0HHmvIJflgPvFANoXTwM5iZNJv6CsQhjaKPfSaClVjElqERg/uo8cvxYu
zlUSA1+iCRS+MrZAfVKWxsRDpB/FYO3BFStoM0PZAGlWvnPzAyCY+wSiLHFHx3kSguYr/F/zNkoL
o69y8Uq8HwscHVuRJ/64U8tMh9PPigWo3YfLGjAMCy/3sEk3Cr0XG8nR8+sACfPA3uKvkQy2Ssjs
6bTE+q3Vd7Z28yXUG6HdYGx5yFGLXJGksibnkli44KSXKVJ/sC+qX1uzuw43syf7Cs0ocz/+35bb
MNwbdObYYDDPQE0c9fVAzYV7bwwemiZeozlpYWqeIqIN8vwIrOvObEjVZ4/YRz0hn0HN68ITOB97
uuaYB5dji1rMrqgK0cNHJ+Be3ybrg0PqpRl9mIiygKM0tO1mZslBy/FGIqdPBKT77/3r8lnLPYy6
F4I33ptxPsg2JCrYy1UfKOzTykaIoRMYVQdQ6XAzQX4LekEcC34SdU8pzxR7E+Wa7l1dTy2WUg0p
xzCzphujWWFPPHgfV0mi0QZlgma+ph9J4M6o1QyMVxOJ/eGdJn0alH1DLCUPCUcBmAejiFMN4zUk
LdPAkRB/ghRWsCbmJVrcNu2VqeRHd0Q9zUbycBVZsML1VgfsOMqG/xOv5ZaH8sh4kWSr8FKvlBix
s5mxxQcJMRLS6Ql9gUocpJbWaPmZlE9/ECCw5TOaiC0JkAIbzdpGXcyBW0EV424iBTXPPWhean3Y
yl8RKAIMwiw145xPVXHENzYg/Se068rSbEf+bmoRlT16+t3ubxd9K8wxtWPmH0/n3RPftyQL0WEK
z3/vEH9VKXMHwo7qM1mnFBJK3Swb42XqoH1h+Fp814NHCwR8jwPxHPCXCJbtRes0nbifyCRcKS0t
CoLozovYGqA8o1+JI6naSf8i/tkneuDH2wXb7HSCI5jN2Zal6FjwXlQnMTtRRXsO0y7OV6Ajv0LM
6g729JrSPWzND2/+Rt1Zo32igf2UE952oIQapm4e5MRbA2t+NeUUHDlWWAq9gN5tf6QPlR/uGzuZ
zI1SbNxCzT8GK/EcK8Kr6hoTxutFZBXMVpraA3WCWeMj0YXao13PV/Dolf5hkH18NcUmY6sImtdz
NSKwVU3VZ3JgbBYbZT+enW3EJ0dG1J+EHs0xyVhJ0jTPJtdzQRHjs6v/IJ4E80FVrrUKFBydGMa8
0+9xDkxIOeO1LVAZZb5h7TZBU3BBm7bKJ2fIIx/DELhmIZNFo5GX3IBD332XfR9uuMn4iAb7pcL4
kbgiWPF+KdYtVlkVxSOR2OPjMrGzty+B+6U3lU26CgCyAhlryI4sS4l+QS3UgOJN87XuMEYN6ado
oAbPfJ3F6+gkdQSkurcQ2pKTrnr+ty86fq5mHslHpoeMOwF9fHIamv6NeYqo6F1NQAeTd5pgCYgR
cZKsL+DvCLhyQurUSUn0UucFNG0eY6wK5xDrMCQbXlqR+FRTu42MAIqgfuhPbORmlc0OlK6ssjvx
gTm/x5T8Or0RJkYc6LmBxEnl5kppaF/hmEw+7zWvNhir64Q3OSy4SsY8Ty8OimG/I1mtl/EdsHSL
feuG8mYvsQnZ1m+LUxYsRlgs+ja9HVRhg/+ACTB1ozYjRfMO6v5siAJ53fr7fWR8CczrPe3UnpwM
6spkF7pUo0BCN9/6pituLSPzd1TUzg8BKsp3EKVEAXnd7XzzxXhiiEgpCDDWJj+C9sieUvGr7P+/
EHD4R73YXiNbdyyTtDFktNS560oUxu2hltkNNPLe4BDN7hdzBSKRp21oKn+URUEeQhPjbtxxxfpU
O0m2oE4qnIMaPytxzeUS1B0Shlb5rHf0wLqHt+kRmwINBRf6R+1cK1cGQBnh95JDiZOIP8HkDrr+
wXXhqbKljZPYL7f0MkciGq8jO94p+IM0qet6Gz2Qc8RwKe8LNp+H92FEL4+KrBOTNf+nRnMNhqN+
ki8XpEUM8sCtGczj9bqPFNE9uJUQx1d8i+R86DAbT1GRdhepR9+RhR+onH/Ne6UGyux6IkIqFzJy
cMNgM2oUo0zNHsgDBVks/+HMR3jsbxjgD5302KaAOoPIV3y1a8AMamcY7GoA8OFU92UIxsNWlqI+
lFiHVj4UY3rN4+g9ICnORU1Jb8zBB2GL+VBDT89BCNJNw+UHYASNv8phOwFfIoLNvjjhDNnnd80l
0boE02loEeDTNJODORYHOaQws4UbhR74LKzZ1vou/aq2/1LQlzGK/RDFTC1la7Bcye6gHCfD5umN
WBHheVOqArN95wuyaymd1E5XuUhpVWtbEd9OSDGUeRkubC7gRqvKBGsa8NiQx45pJEX4Rm9U+1XG
GFFqqLk3NNxBqd2LjYBQXP64mUxhksLxlb6zu2fpsVqvobnCMmEOQK6V4Rgb7EVe+K1eWHlcDDXw
IKLVNXrfO+ZzeLifa4r8MrFPZDGWm08+UVRtGw72+y916/Zdj/d4CU1aFPiH44PdpByl6MTunZLg
PbRlB7RcbmOXbwu3ydThzFLNlz/xycdx79URTyJOya8wAERdJfyA6rIZ/Et8jJpp50UfYb38IW8+
dlVwKcufTgmZRDC9s1FSOrtraz+2DhGSQNyNgnMe/k80LrFGuasjQaKH4iYgEyZ9i2wSc/ZJqDM2
AuI8+7iyevb3bMiMcNSOwAGHZqAQOTxSSQzzh3cfKv6ehtU+V0CCZ/uVwBME3S908+UrXn47DfsN
B+ZJ/9PYDnIvfvA/q5pS4GFxirYFIUrwZf3DFtpolbWvZBhHvsUYvknGmxIjWvCeLnytLFtgrQsB
xGsmI4ivmJA6PyGcP0SjKOxdsKk6Mm2W39pIXhh4zu5SZ+5gwNFV5NN8WsWCePdjkCIy8ZklDtNI
7t7qmxEF7RIMVcTXvCnhShPkyPY0IuRD3Jitt/3JtdzKfO6jG9O5Plh46HDePi/4Pm/JXd9I3IKP
C2R1lbi6LpSF0T1QlDB0Tr7B4ggQUbHebr72ym4z91dZH/EkAeroHmx8U/GwA0VPh+b9uHvIoRAV
ocE/7OOW1VEglLNpTHcnuGTUjb3vZdRwlaG880yUxHEKXnP6K9Pkbd3Ic2PnHACE8ASKC484zr+b
9Z2Hx2FGStqaGsN+pzOKvhTOn1gtUmwGBLPuVzzQtQ3R0sWVA94DTAJMGDvp2KL0fYHmVbxai33C
ogVFZOCNF0N9YHp+wskfS/JtDDi0K7a9F2iDso9gXHD9KT+yf+nv+AdIOCO9iYmtCScoKpe3wEPZ
OeCca4jUCyQXg2bDB/DQ1wOWxYtdeBn4U+N+bTNbM7+yGOuLIM0FiKwLfuLQx6BDGYlDKlUAshto
B3W+b3y6sEJr3wnobIlvQxfHoUTbhji1CWs11RVqew/7kAU7NIlTzbv4B7PJv55XC5/P+3L66UV5
+GYyAeJ17iEb9y5z73mHoEeMtNNUxeF1CoAMGtjGGnPFMVGx53rOgI7KvaeS4CWGium4coP7XH5H
r78Uyhtg2TSd7pisFsY26yoVaT/+YgeDYqwLg4nWtSijYIoycvNyU+MX8gszxDzarODA7bPy2rnT
aIrWVF3VIpWEfeR++voAB8HSkTQIKV2kPSTpRuxjXkffaVR83QGJfbblY0yZqMCxQtmKkIleqP0i
1BKMSNJYa9pMaVKKpQ0my4yvQTx+IvjgAqQ1wKySuwXVLAenGnIm7M7M73qb692Th2Er3yjbLw4L
VarUtlqtj7HoSaJWrYnOMxvCbVLNc7nziHdvoU+1+GrGxMjwFnGt6aHso2meEB7dnh80MXO8n2Q4
ZKsCnb/nV+dpziA+zlFSjjKeR6yO6y8q599NOvr0o3s+Y+UFaZDj0hqza4WlYQ3BVoryhheYhMIa
ZnS/KpkOEFmmU1GzTa5VIA3530FpGzQtqwHyCmTm/cLkyMxZd9LrVHcF++B+yACPRo8SAGEwdg0l
DRQCvm5VzwysKG1OMcodV1YWfK03qUHMnkyQwqO8DzgO4bC5cFbsucGL1Whpm2fUse1qCccLFzoj
/eRnOxS5f7IXbQt3MMzdIGid/1SbvOhIR2d5mBcqfGhlBhekWL9CtDhebhLqUqXhCDsiqSxOjT1i
iyW8uarpuvEsWteogI2QfaLK+gJq6c8IYkChZodRDzmBOVVlGVzFwaCbaeMda9DrneKdcsDXnI5t
kSaqNcEXneH0Ng8bYWIWbqVXTNGY9u8X8Sh4FMZBrDQrIo7CxVX6fsxjuOw+h5C2ZdDv0EXOkO83
ShxA7z3iDY1n2ec9/aYf5C4K4uBX0cic5dIyeJpSyb7hhrj0PQ68omF+9hkmU/p+psovE1ZkDr1w
E6/cMUAmWpCoMEMB3kdFLgwqJIjpZSbfJQbWxUflDDq9sKTujHDB2D/TH6JRuhJcaSktufdddkzp
v4HZpSG5tnCFwLzMqW/7/QAH4MkPXbBbGnNYKg+/wEb0H4l7Bxym1DCbzeNDcw26njtHfeFvElxb
j/qMlQ4lHKScZaAO04wjgYSH77VMxJ+I6+Fu23zV7y1Y7SIdO0rs2VBL1Pbu3xuzhktZXvS9cXOV
LRZgam0NBifa2csDDsgaPp5BnVWiV0nHg5QrtH522bCns+9PoyNPNrs6V1KxCM8gN/bP/paLptxo
jN50Gb0+rijhdGzsVxPFIMQ+p7sfF+qa0JuwTYPFTM8hA8+eQyTKFZComxWzNxhyCs1/w6Nt/70D
d9ZIKJi46M6EhjmkXCf2rwRCtqtNRktuiitimoVe3FZRtC1o/FOOn34JMmMIYkypLO4F653bQb4y
Eyg7xsQAWfkc0T3dtq2l5DzX89VAqeY7AIQNicdQbfd2/69A8QNtckii7ODbkAd9qoLAW7jo3iZX
/QMJ81hBVFAZufS/SeCKOQpNtYFULcY+WdymSw9za6Kqxv4oKj4UMwyDXWZIYNsawWGS2po/Gt1Z
iHoYQk5kGFH7bZ3BKqSTbf28xTlyxVC1wJW9CcRtq4/+Kine7cQgIuzI5v0s3KGARNxpJL/czdET
nIdgv9/OzoTw1cGmZioreTnum50770+tlyGnkFbOLvSMEY8U+IWyX6V3zT4hdJbQ1e6uL9NalXAZ
2i/HPVkogSlBISnh5irhAvWztXinwyyqMkQffYYp28Gl3XkhFRWyS+Rei80Ex+ypzc83OY4tbYT5
4fgxHq6FQW4vZB7jCASLqRA07bK0RCtSF/780HWX8ZiVixpp3H8IHXyLwWdIEfVpRGC2XHo9n+E+
QYFbt4jiiNWTTaR8WpoFcZN2vpyMrdfUTDuko3Gt+XOVRrNf1vIZA3vTiSiKdtZl5MklDt4FAAKj
628gV/MHRFmSHQlxobWsKAccDCMclaautgpf+sw9M753y4UONfxKWU7xXDVQ+JwlBZzHJhvpCIXR
z2oBz+efbA8cn3A81fKocvQv1WWase6vCIdrE5DExrA91T7BnIZCyAoOnLtku2NHwNivEYfF6y66
WSLrof6z3RTtN1k9WN8jTWffPNgtunQV/8P19+eh/96snZv0CDiNDatZHpTA7kCo2bgh5vuOsWBj
DKAy0G/fUXZ0sljpfZ18hmJDXXSCNj5du9JqRXFTym5ZoqCB19kITZAVgeBZR0QdT3sYoWlKN87C
QW1DazH9/vJfLJeChmHNTaalJQl0KVVHsH3U3PTpV05IZb5u96W3VPOboxC4pgUfuAMkbUUIAYx5
6vxNLasE7+Rk8OXKnIM/G+Al6LVbaqLNrgbzgEAiuDchZiOlG+IGz7hWBex0zDg6BmGwHkjv/iTz
p9AoYUdNFrJhpvzMPnQQCkIE4kftafxIVBQr5kHzbcp+Bakz3aH8nMvjjDArydRjgQets3CH0OTp
lwgPALbZyaDZoF95qOnXwFoaqwhWsKK5KsGdXBI/ImxHF/wABVQRxtYhrmijeWcKd6n33zJATzVi
4l5emw6SW0BxTUtpG2F0q0Oq/+4wfTFegUIJ5wRcflVgAzptYOnTcNd/ODapBMiGVKLGbdCoa91j
wEbtaeZWn5cK3lWmi3I/T8cc+n4xWjldS5B6+FC4zotuLLdcqHbIsAqo+pUyX3cJgLZpnW8I0tSe
IZ1ix1o7DssnnO7H6G9RYn75lAquPfRJa8zMPf6YlCvNNecQg3dGOF5owewptz9Hio1DwkBQvPnh
L7dLipW/A2nCSkG9jhoY8cMokAPp3dCpu/93WlXNfNMHI9zhe9JqzfAPka+iNFZMMG0AOlVohoS/
7MdbK9s9NJ8ZAxkT5vjvs6WLcdEJw1YidaY5UYq7IDa25pXJXi4rsR0MPjZEE23xPBkosqBHu37p
cG7Qc0z3eFdGRPeT2YkHJRYLsI7EXiW7gFhXRz3LCSN2f+5P+9nkI8x0yojsi4d7Wg+gxv5+g82H
il48OEUJldrQ0wXSqX76Sjt0QT7vUVrixvTv44OPZFGqVehYqDdFjVDx+uiIhfeKdp+U/j3OoW+z
8BO/XcylhRZH4oSk/agSMdiDBm8UNr/oPxg+SYSYKLZQWkxgpVy+BkTN0yNedomUzW2br94fVE+h
wP8RWrgXzM/xvSJczV9GRNe21CQokYVMHfZDDsI5qbXYWyymArLz+IyJE47AixZnV7qKZHkxMcQJ
6YBwRTwbGaHf4IoJEVFFw9KnqRUTgpc2haB2wYxjYA7PFWj0qWX4eJB5ClP7Hyq5vgUVBC5YEtSf
NGFCj+Kv/JIDMZ0bNO247V2I882XI/R+2W1VzlLQgPCz92+/IXJArCqsGoMBwGOLBKj/gUWiZklo
U1R4Ars0WV+N7JaqNwkSV9Jg/0SqS+5zuFcD+pKCIZJIA8u8uypIpq8GDOlFcsRpbL/Ohmk+QFFz
0FBaflwtEQ+76B/9eowF8dMD99waGaYaD+VD+Ng7hUW9Ttizb3cxtxPwlG17A5H2S4V4LgdeN0eE
oCJS4RwDmrCYjb4/Sj5z6ACwK64liTqlxaeMWGh70cHXxtnULsT3ibIqSuY2GD6ADKtBapwFNj2j
KN80R5WLSAdXATtAjlf139VcENf5JBvMz7tZu4g3LanZ/AfxQoFQeAIzrzASKCm4yF6zeIyks9yL
jfn55oT4N6DI2RC5vCksIkypu4oT9iAzVxLxswFrUrc9EudYjdE2MGEvNrulBmNFFMLgqz5kLDBq
aUw9kwQ+ZBvOaQzeSrJIO4OaQ41eETMupUZz40TxVExPL43vwHXZSFn5hfPxQ4af8WrixPgeo+l9
TO56nLs/Npih2ZGGkzezLS/wz3hwCeP2Uq2zVRglvwkTy9HZHns0pmqcWRvxIrEw54FX2HmepfC6
AYA3DmpwKdbgug9XOk+NLqpxjuqn9SKZb2ISmvbuwfa/zGaZDvc4y6jaf9hVXN5zo9IJS9xZ6um1
c2+qdO3VTEE+YYiigSiD4fpu5hocqCI/2N0z9O1B+V79Trpo1In+OLhLxnATxujXAGlcp4O4ILRm
X6oNLGLUxygVwEGBuqiMIUHwfk/0kKIELtDe8OM4p7YI2TGOfT+Vc64Wh2mJEKOQzaaZdDzGTyhI
ZHFjItiuP1GYBJwgiXmtz4KYem2to3HN+/hAlhQS/gNaFZRIOQ84wS2XHs5tkgJVbI+guM6Ye+UR
V5kob9Bw+P2kWb23zaGsMde1NMk8zzTKJopBE5KF0Kyfr2agRXVq9tGPcEgUZL8kz3ioL/7s53YB
49sHX5eaq8ETPEk4YoKut4m08IKqk3qWLQE2JuDT9Uu12YPglVmVul2Xi4luoGE/Ng2yBMK22MZq
nBDFVrVCLOvFT1hekQyOWQuuxXeIXWyayc8o24hZSV6kz4fvK21eYF3HSU6F9i1cLdoIjn9fqkGa
ng8GIOHSU3W5o0t3+ckgovJRbYj3nghf+GND6ueTdvyzvEQYBGyCj/2z363IW8joPxsS3lcv9aqA
04ft99+CzrYefZveTGUHtn4mraU60A4s73DTtptA0jAbFDOcKAcogVYI0FhLWhpgkzBDYzE+jDFi
eOTuLehYnVr92FWQ+owjo45xKNSRthVT/XN+xTcEZ4AUp4iYqVRg+7JbaUjHsBVTr4cs3WQmeUSu
PgpOSPCruM67HQNSQEcjUQSzKeu017HHYoADrzxadkthY0A57zNOvX+5UBpL787gbpZV/YwWKIaA
nW0ludwD7vPPN8oPiiUyv4Cc6t5SMfALqZrTjJWu/TATJ2Y0aIEhXlpcAZ3nYTwrIpPmBd9WgpIv
/cdmfFhiZCbQRYDZfnHyTJZTwboWJ39L5+4aJrQCxTv1vLY4TORiuH9uAJxmkczL/QpMjEBogWuY
0du+LVWJvr+a+wDErxWjnGVKJGkd7363j8Wm1t36dMkrCb2Rd8/kEyrWpgV8ZAOHSEey4ze6bHRC
ukdxl6POOmUQ4KLfpDdbcgpXi9DILU9qu8UE1QL1RNj5GFZ/KhhhbjOdWoCwDy+bveiE1fAfeEn8
1m1JdNrR3S1I0ehqLAbxBvLnx4XDPnMiP/KM5oyPyZPCIVlR7VkhkFFSJlir2FwE9KfdrvWlPukX
liIrVh7/K3ucNrINJgf5V2pau750x98mMz9io1fLOer8qG0YiprHqPNPT8vwd+Skc1NfCydsvU+l
azPW3V86FaAPMaxgrUDIdedyXnJqegwT/acLUVGc6jRkEWovxUb2wlSW7XkrovtSpngVlhp7CiUq
OEuGS3kLFqJ0glX8N0IhTlstvDmE4AmKSV3IXf5t2+bKCbjqKcRQAeOvXTQmZGZEI4lBW1cqE2df
DLU6sta6LvY2JF7LF9Me3fbJDkRRU5+AHAlXKSZNu2CMqPPJiZHqw7ZE4t+4Y+0umYF6c4YGGMx4
09p7XxCrKLkPQr7i7U0xdIAbhi6f7zaa7mVr17oFrcNHe0le+Im3rOjwIEh1mT2NGAM3uTu1sAnl
z35ERmIe+9/uITHLn4DOR6biiWHVtfCoUzqxcX30oMZyfucdETdxtNwcWN1G06A4uW2V3EFjEGlB
tp4X1S1Khk+J/Bnp5ywjHaWypDEOheOE56dfu1EjoTgKNQg/6isOQvlHftV0dc3ctFEb6gqrF+on
plbH2nKAujnk1vweYFySSGeMpSuhCtnYVYkjPd6ZhtHBGpLGN2bQTKm4kT/Ap+jwY/I6OEXv6kos
n+P0Gh/L5mVU23ZhgwORUNhs+iemTXy9ywdniS+9Pc3bnpNBJ7SroG5BdheVZGluLTdCLkV6y01M
M/Y8vSY4vv67zj0Ccg100i8tkoHXf+4Cfq8KqFG6IWeUJmaSgKSB3YJferECZtVNNugbZevZMYgG
LJMtlDkZE2FPbQxpPRHajAqO8Mzg13+UMRqJYbcFZQQ1lnJrMBzU30ezW/wuM2vNcqVUgR+UECEZ
0Pun4E8K7T4QCiEMnR83f9+QMIFTDHcUl8+Zh6ac8OXusl+eh1MlG2chWMZhVkQaLW36VcLi4LYk
25ICwkjBnu0kHB+gs4p6ZEsjX3rJgJ2mUwhrxw7qSM15W7fUf/fEDS9zkd1ePb5Nk6u1bMjzeyks
EDUJFuTgj3BSY07vj8F6jssQMppE9aIJnVo0aXkw7yYzhZvm46dEcGF2RauQY5sAcTIhZzVzm06t
F+e2thQimheMDvJWcNMcCBViAeBC6wAperyP+icgbchFiwha457Q/wnsk9KiyGQiquzWOz26qtVA
uetqQfzjd2qsWdt1CU34HZxDCzH059jBBvMGftoZWZgzzc08UP9drBBhYAZ1wjfgmG+BRsEBDgdu
zPiCWNEgZlaG7YynoIMpyjkDB34iO6o6eTi6yQdO5LgtCFEGE2vmlY5Wlm/Z095FElYXTODaLGmm
YD/YVUY0ExCJ5FwZcFEQOeb68seefSquFB+fxQNvO9hUppfeoDjVGjMUawDycKIY0xqP4B5nrQGt
rNpBILwf1rGD+vgVXVFt45pwZ8dMN+QpHXcwXv/Elyp3Bo/3te2f5Y8Q0+NE3vpbb/mY8E4MkGL8
z7AiAmvV0Q3MWkIXliPHNXiEDJhk29b4zs8DN1d6dqBNoZ5BeNzM93isYEAiBdbQvahVxp1DCInB
YesMwnP59DfTWCSsarAIZysDkzSdHql47cASanWnn25drPlsnX93yon/kXBGkIwr5WV1zG7M7Si5
hMibx0e/VIbGbDrnS5r4L2cONC2ncl8lzbNquetRKqwmSnmWXbvAVrl25VZCXIV9TtnYRXx6FFBO
N9pSO1HX9lEAE+nad/Mo75uJcBlkSYIPJldhb3elaN8AdowD6LMvKGYzGhvVPabbSnAaU+L68BAZ
sLcKp2dwaoPc7o+874t9JW82W13I6+el7iYvswl8sDEtetf4uS7JSY51ILAJpWie+j8O/4NJ205u
WL4IVBVh8U3pQM2gDidMj5f/D0VyEF2EnjpzZR11v6v1BGKHhkNdtVGTwqu4e2AJWSpX/dlZ+SJj
3BiYXY38funEjfdTERpHTWLWUFAWtz/m8RCFd+E96dKKRBtpT/aaHSntQlut4NU074aKmJ+KVLF8
sYxsocOk+PI8rPa781lld5+dewiEUCnKHi4FWatM3Dajd5aQ3SNb0UvahT7DPYnJuXPHSgDqeKxx
dzH6olCYo9WDgskGoVYNDYFWzCSBtNEFvJdHeytdQaMLn0aYXZHL8gvYC7Ls+cb5KUJkCcWPwzpM
KNAcGbCoLGD7rV/9YDn9oPjxCF4epvJP3Ee8Y8pKcIJunjVYgFyCqahIuAvuIfm6NJg9at1IrPfA
206BP7htZbTY+yAtlZL9o9Xk0KZvi0GPmbf2ywWeAj8Q8wrLl5aNOiXESvqR6P91VFjvo6LqsH4v
bT2TYluLX66ACaWeeCxmZDlqC5ziERRA8LimsSnoLh62NiXGiOfgb/xittW6+akGwly/0yyqW4M2
VjODc5SB08ZQ9zvuf4xfMRnOD54VxUWd4Kt4/uZ0TA9h3/y8oZqGQzVEgqSMeMH6I+OM2ZstmeXS
CzcWcRTk7RphaFaQvrQWyMEHDUkek3Uvt40Yse8fEPQdpZLJ7Ho/JueTPUphDbsv/U7D3/RBwoe/
/VxgBpTsjTh7i7EUXSoe22BTxI2UF+V3JSUIJcg4ChjtxaoYq0NicoDvpZQlaV86vidoCLjtX++2
CWY38RXldmhJhwBVViqk8Vqqia9O7MPJe5yujimyTQQAiRHoTTpz8E43Skn53ZF0Ujy0OSJmApiQ
NDWdQvi2gBFY6TE17kG3T6ert1lajWvXPGmFgczqF0GLHsPL3EfcNprsTsYHyOMO+ZMGFhLoVhoe
TTB0dKYQrSFRGlM6RKMGxA/Ci0Vj6LTMDM28YfRp2skqL0UyoQqBno8+nxFQqSTg8xdghA/cI0Sl
ugmylYjwEMv/FgX2QV0TPCbAePltE0i3mtfAscfaY9nZj4o6JAlqQg5MiGBZ7Jw12/UuxlNSeWNw
wUuuWCcjYJC0TYEpmnpLjgeSd+cRF6LD0tiOH6gq7Itvj0jZCf9R5m3ZxvhOIsdhIbU9Rbz6mN2T
AoWBDIbbmSP10izEoX09jkcbwdeyEcIL5Wzax9wiJtrP3bJ6B12LAlGqltK5HEdBD85RQCMuaDv3
PAg61pCCoi6fzOCysmwHp+Kxm9wpuhKpxdLgM1OThcBhxI8FQZ7FWnw46WXlDPqmMJyGCzVNVm5W
XanR7Y7ZETUs1VQbab9CMlt63vPS39ufIaV4WmEvVYKewRExvwLJ3+Kcni6NWdVbpCsulRVD76SF
bVlCULHjkDiXHhtArTs5w5N2Jcw6IFvmRDGUNqDaBq8cK6BJV+dkcwg3JXjS9zE34NXDjgeimyN/
fiLko7cu4Fq7QMz61Hemts6YtKvtZ5HIJ0bpRH0hxzb8+7h0j9xfuwGQ5hi8Ef9ozkEk6tLPImCQ
YEnYYDmZ2gJ6KHD6eLfKxuhAB57+McqHO19yntJAE4V8mY+zpe1tGs9BqxKvSlpRDimsZItafxFB
LmZuuYW+QynAOeUv22G1KCVYx2ctpkFHNZSMz7R9XW3euV1V+pVNZcA3C9SS5IwfrHDVZvGWEzNH
aEtKEICKRo76z5pUce/WFKb3UvHKRSY+v7qvh2nveV/UXX9osNz/T0M65mw+qgVm4EO3LkJBUsOt
eMLaty9NdlsqeMEqCDaV0+nyTOoycFJ0GiuQfnk7CjgkA8TBhI83ZXYoAFaRUkTBCCohGVobGEUM
qwfD3kNa15sDd5afIDLRF+TUgELdQe43+bin6IjkzCWqOu/DI8hoaMzqWNInFV87iKhE+Xi3rjOe
s6fpA80na8l4qvNXmm/LZVKYhW5SspACntCTs9zSSgOLcq5RZwO6No9jBDC5nI8AjjMGjzoZwoZl
A1LBlJsjMSBEwJRHDEsiVgwjRXFY5gpIPj472snR4Qh4vaeWnjQKH420Y/cvjpds+qLbPXCEYUhf
jOW4XliczJIhOBMQUojAnOq+SA1chjHveWRrBBpu5XH6BzmZkzYQrv7aPfFnhk0QCOp8PKdLosEs
viFHj5yTLIsy1EMmSZnU+An+y7HXJuS85E2ztpIhpXTk6Ya+g5cC/hpUa8JQYvxUXOOEmF5fAmg2
PC6wJy9vErY9nPTTC/9cSoN//qr1Sfi7VPEjVjr3asyPDEbDjbdDMxxNMfZA3+0lrJoi9Ly3NcQb
CKbQ1XIkoexnYw+VcOu+saVGxoV7oSvWTGTQWeTDPvjOBtS5BsfRipa5jKb9cPIXdELBzP5Z95Qf
T2lZShkIs2d/cfQ9k8Y6RyqHwFJ9Gd9tPHdA2ye3r4RTRI1kA3sIR8/6W/3mGLiohylAFtC6M6Mp
TMWvLfYStBDGtH/QAxPgYWvOHHi3QUKjK0ccHykNSdCjG/I2jEHLMCeFaFaWdtG82cC8bgMVsGVX
kN/XgZ/UMSOI3fXPXnY2dA2tlfIpzKXcXLiDhJCKGrgidXQ6HEVBZrJmiMeV4iUzVHx1NZghNqDp
qEzU7khMy5KJey1TPUYRYfGkC9dWI8CEBHUgZ1UbP6jzuhFh/gL6TP8Di1zFttnC25TaohzFfqzD
5/x7f9kHx/gTEIfoZ3t6BuzvzzttGEIUubc3QTrDJrLd7ViAjjzsbxox/jXdvqwqqhl+vG/eFo7M
Zy3UQkt9BFGsodWQK5R71HTFP46fq3NfQSjpKW6PMOcJArZM0Qn31WMZRQjIXAAhQnGXHwBLHmY3
Y8xKWz4/SRNJE+2Zmk99LpCRgoKYksuW2EttTyaEsRO9ldWPd7vj4I0Xi4upg6yGzDlKgZJTKj6i
VG/CqlSKj08rJqRU15XCm/Qsgfex4fxBhbPwbeDZ2un0ojeG2wiMcleFJ5P+5gyvGOIKkscJe4L7
rsIhU2fdgYbxQyiw+drBZVnM0mbxbCp3jSqfkYzdGfbRTNB1o0pGxbU34PU0H/Stg1AV286B1ABb
39F9LeaRmYdJxleOAaejNhVWdL5wsbBIhwXFo1KWNg+AOVbz1wNHYsxEtmxl1H52YcM8dJMXJSur
7tn2Zvm5ebe1HOmbVKmz7H/qczqijRGfobr0a7B7asLq+nQEDpxAcwR+GwlfwDbA8QEkMi4iXgao
rMzJ8oFerlzahZtNTIZM5ABBEzsbqsrQrPiyf8O1XyITHna/1/3jd1hm/EwYkFPNrxTwsfKQSN0x
eH9QuH8pdGH59bkyHum3uYUww0o2iCPbYvhCrs7APYiXJchNT6+p7N7HJtZpvYs/L9GoGdghoMjB
6UYTpiAUXdR6m6lsukXLjcUJ2v/ARYKaJjBvQXStGfn+w0V+YNhCWa9HIHZQEFFv1u2iPGIAGdDm
ggWy/S6wSCFlvexGvsD4u/2Ty/MmxHod+vkVH1DkHixuPSaRkhtTJavqlcG/RqPtOvAPl6iZss00
Ni28joatDB3TnaTkgYf8kg86tWoprE1Dp6g1SfiKJldUulM4dYAhgbck7i3I1jHys2vmQy/WTjr3
Db5IBO1UYNktMGFRT2qvqu+GmhEMSuIyzX2ibWZ7DYrmsLTiY7qaGn6/qjeJrqN7cVVw+1p8v/nR
3LHClQWqPRzE6k52TjD1iDD1mn03wU6D1182lE7ghQ2RChEj7hz8ED6mrBDdzpQg2I2d/oNBbo6i
RgPWYP6WOys6A816U/9EKwRZfkVCeZvNdc+btvsvxHlu/XKd5VYlz1vkheL52DXxaKc9fbN1svFm
Rw5Kj04oQnXfQWJc+WG4mSDBs2Bnx8tLW00QYke+NL21oZxZ0iQpQ5KqIQlXU5544HJ95DN1h5ZN
EAShXV7HW+NZP4BtthcoTAm2SCLBCEf1NbGKz5nqu76hOFS2EKaWwKjx6zQRyOF2ytVKIxB0dyXO
BVT4C3I7QRHQPDv2vINJNqqis/lhIhtss+KvxFridlIkuDrqgWD+W7VwEDC/NM0JEemCeYhVuMhW
3lTCyplmnugqSgeAihrcqmKUL9jdBxwziUHnqJUMmfdy297ognkGqn6mAM3Vdvhko10FE5S6JzMD
h4lRGpC4PtFelgwNTFIWuhzVb9NrdH7KD1mFJsNnAokavTdHuGqBUdLq8db+vt6xf+83X3G2kBFE
sloQ3kPlLs9lhvT1juJrcn5I4yjwncnpGL/WapXmstPb0vU5sC2vN2FdK/xvDXQbv7GPMm9OSF0C
56njv8p6QqErMbgfo1w8gWYMV1c7Xev79c5BU4OETq+3x04ugkpj947aiAyAP9E6OOPQTsoo70P5
Br3CYc85S8/BC5X4esa42uEhiTfNzP5Qt1pXNcMpjWsoNCsT5dD4qXSWbc7U+eqpduwFYwzI7vPm
1yq2Pnu+MLDdEh5UVdfhRmVW8uQOhE7vmSeO5UwJTJgqZo+yAAl91DgHZSpw+za/H9FZN2sEwQju
4/GYk133LZSB/a21Fei3TY7gGVo9wwf/c8vie+GxfuAOD3c+qqmNwOaOwe+1pR23zpZi7m+Mi6Bg
lJVml/n/N9TODqaZnSIi8OlfSnBwoUVBFw4CPn0JIGY+ZR9Cykd86m96Q7XfXA41cOD+b3VJHgFb
SPgBg9Nng8vZ7dcuaQHZS/+8lHEA+RnanbKW1o0DB+T1vO00nrkLLDDUAMdL6LvmdHtSmHO+oKtM
lJvcLyyfwDraYp+vU9gXbdAILXhfyOBkyjAiECNmh/q34ptp78VNJyHhxurI90y2XyWZraRTYeId
Lnj/K75k4b5tH6aUSWVYHR/LzhF3ipZoJ7ceOhF5lI46nq7pNybTu8ECI2btRXzE7rC/az8iki1U
QCNAllp25cB4BtmTGS/aYBYdKI3JXyQbQL0uXam+7TED2lkdgWqOBzGWXE5NH/538FJXbDUk4jZm
UnoUWHkSVTtYHy4N5Z4Vp6+CHwvHG2Zw6+53Rs5cmLIhmr9REhUTKCRut7MOqR4u8PyJdULz04yk
MOLhWAfPZUaPopWrZWeKZ4O54Xm6wDv9PiwQLsrA78G0RDqwQ+JAxWnDPGT1GD06QXgirqLDyk76
f2MZxtrrEQuqnnxR4xI+/VeXVkwPtIhVLQgHBSB5iiKE4Wq6HBsr6wPge+h0H1gpKRGBrG6ELdXo
Za7nTgmdzSx5UmRxFfyfb72oICWOD4oYY+OeHTaldU3fT35lZPN1luxjYRAwi5ZWwiJcNkSkTWq7
LQ1z5fj4x1pPQR2vBmRUDA0TfLcVLej9uwO2Q2GsW41WCFdFYnB/5x0tXekXKB2Pno5WVbr42aQo
3G7vosaqfy2Oz+ACf+820rg3S0JKsEcIi6RgQydiJKzeNUg4s4jihHEYh57dxPflRoJqLDWM0Y9O
Hbx4PsRVvspkole2fHb/nUj9kk4vJZZ8XVnkUWymkdYjeRNoObgsQk6Ng4eCJeOLxCj1A0ZHhaVA
LeWXg3ypvo/DIwgt2TQ06JC1Nf3HoSiYk/bJlfY8ruzNdh2m1jX5+g9CD9zgeN9IKg6UsDMOSNDp
cXSarujwCyJI86KjF8AVPPUSo1LGwgbQpSy1qbAx04h0YqGNZGNqeTuneFfGWB4hZGFc4q4qtdLc
qg7SFnz22A/2sO7xanKlCaBizFc+Fh5ki1JmC4NYSPZfMdZkhpuBMFnG03dqOIYVYRdWICck3bZq
7eAtqTXRgnYsI8JGleGJM4U2EAFmHzASnBjtq9rdXjOMhB8AM5EPq91PlXMM5WzVdwxMB+yrrLZp
QFqfc2Sup88g+c3s9YMsygsWvWdN9as3mQmRXZp3FKZy74x9HOXa/sNA8Yut43zpWr41WKzwkCKQ
UykPYxxV8csdwG1pEvaQBugAAwxhnEmJjcr9BjIzLgFgqXTHmN/bHLcvXQt0wtN5ZSFzfSvL69sn
xCmjCxXa9iyylsxvwQLFSQ3SULNzgYhO3gEc1ByEhX8cLXGLK/EFRfjAl4yWPYja0QrZ53s30kPu
x5Mpt/BOv+cq6hql55SBQVeNwJhHfhXmRQpm0/WZ403dCNLjlU7TKF5SObumec44d+D+1hyIlJBu
76fJ8XN7XLKbPH15akY3xkPKq+M1AcBsTCf4LiTTZTUxkYaNfmG9Bd2MF7Xqb9XDmVKgetzYEZiZ
6eAAB5Cy22j0f1uVs06j9IHC1vfmyFuriSrOXsQ/SMTVXXWuMfWQryibnfi1A3PzZ/I0JKoLDEJm
WEcs7Bilp7urU5XL/yDPKcK05qcJR94hBE8hFHkSyTZB/D6jZuem1d4mssjiyYVCK8Kly7HmTTyY
jKK5OsiKxdvcq6V1k31KBSa743r89kERXrMK4Wffs/CaONyJl8gNhVSazBzVFSlI7Vhz75Tluxhj
ZTnmpM5A7edaz2L3/5iMuNQpnH0Kjzzm0GeRY/wHVIIpDRBvfQ4y+sRgfqG+fKZcmqXcI5sNqOCc
cb8uH0Jlt5jM4ED/2OO/T7UtqMoniOjm8fkbSQQCcCwcLnw7ZeHydLFswhqi6s7Y0JtT8+dbHtdV
+Q74U+THPUx31G4G2xYEqUdVcFQkAiKorlL4LDF1rD2326KD7zKW1rfbOArS3u4OrHFpi+5BSifW
jMWlm1Fk6gJh0RT1ntI3uZqS5Q5Cy8jxK1k2OSk32zWqwfKJeM6XEtwTjg5Bh2VZfP9VvduJeeLq
Oh7/RL5BeLSXSjbOx1+hO904csLjytfJ43ctkcqv+pM8GmlAaQ09UwbNdPVScJtW+GvCLC5Prn7p
MMgVwJW7hjGxDIHt+7J9Y0nj6v/fe4SMoT4XHXpWGJDrZ5WYco1KMT9cGxis2nIcKuySLxt/Ha1b
vHmBmrOV/dSwVHmSpku+c2wMlhfCWidZWkI2IHigfhywp783bwjZOXu2EQFXgiTJeHX+Ma8yTkIH
V+1+1G8bPk83vzbQk4rh4UGBiOb+Cb+4Gn21krP8ZuuMzlSN3kWOGbbSIfAKggdHWmkJ56mhXbV7
+me2B4EQycJqzjKZHUmj1W4MBEhM8t/AA7z1HtQZ0hN8BaTpPOpC7vIA0sz/W54zpjKI6vosYGPw
bnAl3RLA+QS9R+qr3GkTm6ILwdUa9kwP7l97/lZpkegneUhIvcPDW7mpPLYjFYilaSe38O55HQYF
I614ioHGYlCMfvvSpRmwRW6TP8HnL7xeQo0lZ2QQ4nI5u+p4JVn/jIRLA2i430BrKhYoikD+hhWJ
LA58QkXv/7Jj9FxY+qDG2uZHqpXqdRonq+LbMeH8B9wLbUkahO/v9EsMfb4vb5+Nrt7UXpyTwYpp
XLZauxV1jOLA6ZbvGI8u6+pASwoDGGTdqIbwXAYlqZFI67NiH+43M0/dfHA5Vq2Yp/b6DURSBG8m
YtvM4MVcrENeEBSnmUjxeGjbVVQpL/cDkgErtQ+zQxnGYOxVCdtr84pzPqEHNaXdDplYxk4S3zRW
RQtqzC+7B9h4CAsheB1sE1UmoFKL+ChIgahnp+bRnUyxFaIiTaSRtEX79Lj9pSP7sauQ5bYDsEww
Ohqse1mDIbJvw6wZMeknauX2+vGWx2z859WsIwfBpUnC7VxYC2ILEl6KzA6aVkIr3To7l/L8cWlm
JABBSVDWiTC3fJznsZByVq0LH6tGWqDuhT81YmEtuq7dXUeG2di+0O74ChqIu+WpvL2w3w12WSMt
jn+4JOxHcIb0KOO6sdqchsXcUWmrHhpWZ4a4iATBWERSPwXBGtb7ilpPWkZ857iNEctziUZ1gJ9h
j37P9stuIAoi3H31rUTLf9z8bxvxmmawZyiF1HuTruYANcPTGAsYSU17Q9Y4AuDrq9liQbV563NV
nbSSOjsz58zwh0HNs9mFKHIW965AUYnaDXIXAmHFXe5FFsDTUDH2ih8xZjVVMLT+JpRujQqVsSFC
3aLEtLyppoT2xXe+sBuoC4l2Hyvkqd2VvEybOeGcVyg8W7xVZOZojoJVAp3WUkUFXTZtLqoIIavR
+tpoYt/M1qYTj/a/1jwjw5vZjM0gWHyjCiMVMdPhXh2knJNC/Ur0RdFd9xJPkar2+sHuz/XCZ2j6
QIZs0Q2WqMJHJ8OFeHQNDjKi4TMtw4VmPy7ZXhJyvxEnyhPtfLUbkWAkNHSSWYHSFJCZVQ3ltuIq
udMjYQiyck0xKlAimugI+FORFy6JT5XhxUXdb2WixilHnPHybLnLw1RrcRmwOslhasJXl+2bu40R
Ckui78k/CjfpGcsWGFH4cyUeRi9q+6xRd//YeSjGv9iETXTSVTrGAmFJyXuYEUAHV2PwhSPEhUn1
U5j9AxsJMhksGCgKhLEDDhqiJQCFrndd+72mkjpi5hlIFJWVHU3hbxBk1TtkdvFcZPHuSZhhHKj5
RcBBSKbs5LmA74KBOQaU5Gp/k+dZRo5ouRD8aQWHASrNUAMLVz2tlPR+WFo90oBgZlnYMGtT0sMz
aU5CBP7ZJh3/mYtYaUGbd3/pEhx1LMIpBHacWiTeUbRHjAvydePz0XFr5/HEmHiuaI/ejFSosUhS
YRHW4VNhEDTvybXc5j/jSpPEYK8qK0IgbacveSIYPfgWCUEmTE+ldpY+oeUxkEg6hyB1/vyyXAvB
POsEaeZADwYDHqXbObFtzv7o5haHGCN6N0i44i9gdPt/acN9DQufL6cKzOj23K4P8HV2jIO2YeOk
XD84qsmqzzK1PV5tlgHssVeOAcJoJwp2ItgsnUyO1QDzqAjKhhs7fQg2OL82YtwZ9oHGwd+jYdZZ
3DasjADLIdrmYMLMOLr79+6vx3XEamPlJqt0AjpctSNtyuHYEhbdJkKR/c3FXfJExX+vOnJ8hOoJ
G9J3G3R3mYiE5Xi1FaWJY9FqbtEJWZnyYaMtkqjzDbjll3BkTFp6A4ILIGuVEnCOJPy73VHC1t8u
W6UVxwxcVG8WC/xWiEL4zJyApI0O1dIFB54nBs7KN31wub6b2DUO7ce1Tech8qcROA9tQ0BVeXQx
lf/T2pvE4Mu9xtpPrj5+bQlEuxye1GkNKZuG7nvLyFs+yl+55CbLzuH4DPXYSodwPawhMGTCwBAx
8liTvMMc4LI8YUQCch8IBB7YBgWNy/5zY05DT5M4ZO0j0TxLYiAk7eDEZGoFDLskmTfvEaCBG6gm
HW47CzXh5hhbgEaMNncbixOOXnqfQwtnDEyoY2cLFXEWJXKUOgH26La4ci0TKijCVzkZczcHiL9F
XvoaCm4ssDt0OeR2irf6UO+69UrRYZCoSyWhX+jPgrE5olPi3cB8k/K/J9e7gW2UbabvDK/R8AZW
azdxq0gk7ndUjLoLzrOjdpSBFTw0yLhautwQcZVfmf3AWTqCRN1PYIMeh47H7WrVifAraKKxe1vw
cMsKIXFncAP0336Kdo1ms+wHYq7ND3NRDnzkWaDH+PQ91UWjJnPBpSUkC19ecdtW/amRp2Yo50l0
pxQbLOMjx683VfBhSLGY0YAgili5vU1CN0/7UbeveYBhasNrHOSM5PrZjVpbtEEPk9N4waGFV/sj
gMImpTfcmONA/p4cgWyuIsT5vuu0Reu42Ht9utWx4n9Y00U/BXvcfNy1Cn86T5w9b+42HQsQwlK9
TE+sFPeU/rSiV3E+XsyOpFDtfo+d6/VTA8yhvh/WEEOgZxRuiOsGDdAuOB2AmUI7H02Xtg39Dw/G
rDwPKkiJzizb8++GK7K4Y4dfzhvtdw06A+8KTJC0+PdW6c5E59U1Fi4brWysFYPtQapKvMTR9fQ7
NOIH55hndIyIgJkRMxJ5p73eOaHq08xgB4BiUWuKIU43BUdcQcKJpNcNsk303kcVe0iVV08pmtzq
EEkdt3xReutV/+dCf5286ets27dgl4cBf8a2J68waj2ZpOGW4AdUrFNqpRxaIdYmr2V7J5BcK64o
oQHwlCHnDT5czOaKk/DjKJb2AabHL91jWTNb/cIlhtuys427wHMXk20UFUh3zzQMD0vjM9JXZKwE
F9wYw/SES+T942NzMGJZtv6nwrfNNWqdztvKbfcVG9nnmSnSp+KZZxnbn6N2addK4sVOiIznD1Se
F+mQSRNN3so+D71qFgjr0ae71C85787fUwOdLaeYRQYWK0m9e6/BQAVi7NOi9FYbGI+lKukbR03i
LkvwbAmtLzXBWrGbyRvZwyLYJB1WeN6QIzH4ACU5TVZX0CFAke97+z5nvlZlJootNu2X2HTqAFyL
WhvfhME+9pNakC3KY0u2hnTurBtm2H1e8t00mA05j6ETa+gs1PlQa+EvEIN8ivavp7K+eswyOWcz
He/p2BlMa03dzAPrydW4STpJJyWk98Tv6I/CS52A6fZAIJgK+0DEjT/2l/cJe5L0MkpFYOGhuI8r
wx0r/RnrtUp2YSSr288L/jrOntmU6Gwvpr8EoBzrehluLUClUrUf3dseNyi0nEM7PPYt4qZKcVTx
KeArUerFowViROe4yY2HQKO6HQ6b3w0NNF2Uw86xiGF+6rk70f0KDZYqsP9TtGNsfUPTFpKUfrnq
Lt+3bPUwicEBKJ9JfubKPgJ9r9TFqa4N9xXx8ntbPXtoklHWDoi6sp1cNJ8HMHJDCkR6eYx6v3Yx
NhBZlWmQ8Y3NgX/bx9eIRM/ga+71SPaHEDMRHRBSwbck0RL2Ib7P9pSfrQM5XB0qdcCzf0rPPlgq
Kd1/QeA6KVr5DTvy9R4T5afix5H8PMj6VzdNjU28ZRh7JYFFlShnyE7eHMFQx3bzLQybDaOAt/lK
43Fka1rpQYdbjsmKtPqCvBYT8hCwIW6CJQb3faO0+v89oN0o62ZWND0dgdHIborxbdsTgBe/g2Fu
dNcJZC+N71oBjVkY/keXyk6Bak/PtcUbmgxvRpWdmuVQ+QZ2VlVnjrgz9M7S+Yk34Bs3ifihzSxB
zQoy0jngGIscj2KlpIOdo7swgEbdjFcs4hcj6TQYVgvR+3WaWRc/5hSb9QyAVPUhahzx7hLWPWrg
lmCE5s43Ax1w3QMR/G3ZucOr87Y+a4tSWKOY5AJoRdWbZpIOa+hI3mkLEJkYZ07Ps2qzcFjHrc04
e2lfpMpnuj3KW7zlh0qo/4zLlA7p6Q/BO+q7n020yDdHr0TWijlzYPXTbo2dFTtJwEEWzPeYFZEy
AFwHudY8Ov4jvL5s897pdD1nJ+B8Ob6KU9dTFTyBR+LVpNXsfSkDxW1RLmO1FrpeHYo4ZdKno3kZ
qxwkJn2Ogt226IGSpocFuKnrepqrlBkqXvPyXyr7Bg6F//CFzfXy45BavDpo9wODTrhw7pmuSqlH
o6i31LPsijy8c9SNHmE63mNcfhhYj/YoDz0I+2YR+TIs7i5LRNh/k27wq1lgw7Q3D5VbsCxllPHZ
fVXixjO/eg6g9q2q0Liy7DR/7soOCtatNBz9/MD98sYIxBFA4STAhh+uXcAc7ssah2VugBEp0atm
2jpmOXXCuWMhVGSPTwFsLZjT8OaKRLmYolgIJzqEIxL5lOxpAPvMoDAT52fHyptBdxlVxdx/F4Xi
bFhKO8apf7qQGk/Eo+IOR2GZTadgiEaiHPuttuootCSZiYxZngkoT27ZBS7VLjcUxmDQ/I8NkZp0
BInoTX9FHeI6gnI4vxwamFzzsuFbwvQZLpiHsc+dTMXftInv2uXo1P7I314OCgspuYzGR+2GxPQ7
dK1e2UYtWrYn/mPNp8JNiFPcnBlaRCAYpwPiP/5WT1tjD3Iw/09fLFJk53nZ7pBh0SJhSfrx1uSP
4goovnGc11oWjKJkwLvaGSPrhjaVNMnWXiXtXkHdKhr/NxenYjSib5jUgL9HbeAPMAK3c4u/3RAr
p35Dyj8nV/DHihw5r/n/UexdyOLdHlF5/G+C+pkUxWUFKdwfUxEZqyMrpOnrsHs3VWgyneyK5S5M
UIRbFC7PvIPCRtCiDixMkGEDHhwiwMN6drZpm0yw4vJpI/VDFlvA1WXYjUX960DA1Duw5s0u1snW
nztHE1dB3jSJ3d75QnSm3rSoQrf7yN/j01ptBdJtvqFiEehK/bnocfc1IP7AvfzWC1LiHbhmzGii
5bn8i0xQBWTY5CjTmO/SWXDZP2xuuvYsSNeqMmDMrI9a9toA65UMEvbA/NtXB/dpXnFbtVg1JSQo
1OI9UXnJ4WR/jsgLL19KlLtbrFaCwnQdvrhKuJ+xPikzrBmcAUJJOE22sD+7/7lAFQMOnC6J8Y5q
5quRRtykjkoYBioy5TzYVapLft/vCMrBnYdBFsmTnKCwqtXXyPYnLNHgFp4OQFAEpNiLb9cAthhS
tX4Ixe9J7SJ1NDjS0U6Lbek132dBKdxo7o19if9X0SWVWgJOh5zcRTJVt5o6Izv83Pjdvq551Zhi
LInoQNm8y+5zbvFfxNNdatNJWvsZAfg90YTr7YUiHDxeavkjX2aq3t4nczGF6WT0XpyjZqN1eGzi
RJWj2BC0kta9PrCwbhzue+vYiCKrHUjkcGu8xnH+SdmjLvl55G07bt+5hSdJAvB1PMctJvErk/Ow
dvXptkSPmagIObUBzdKvG5Z3Bc+tH0z52yk6cz7zffUbN3eYWah7EBxcYvi3n/dYXNTiaw8zFb/A
nGHYggfDZhqh2AfqsUYGcZ6khnYRziy/8tK688S9wGgFhSIa4SMJfzaSOf4BO/UwaWZNfsTCmb/X
H5fzWw8yzEbK6MHUPtetTjlcWUcKU1MjiA+3m0TA92/tNJsqM5t0TsFnd0nD2RFc3b/QoinutrX8
69Q6PBBGl1XfDpJTlwqsiOafmsJO1fVE6kea1BmVBcJdFiomO7C1Imonudx829hU2lkF6hADqYF8
PVorczkxUi4xFHvr7teBtp08wUJeu2hywOdAAYpVSPA94E7WNOszaGs9bT5rcvUqnCsMTDvtXCPt
bGkfuUIEysrKk80FICdnG8p40LvxUwanMqXHP3A3mfqFH0RkMEQJEOJsdUMD/V0JZaYdtNTq+Rkc
BA9PBntqnYeeZ2Rd1HHsLJEPG3FEZpjk2e2LY08LAFLvcFJpazNs1fzmUje/jl3KZbbOT5thiy8u
ANCSboNH4DR5PeG2+WmWpgA3vwiZPunvR8lfuZjdBdar+FezEB40SLo/BLo7v+G8/H1ZBNcjNFQy
fdNSnnfzB0oI4uEaSGn3URWcJPlGRdWwB4IKmnvnkp/X/8AdkoJnuJnShG1ddmlv9380xamUbMHq
TvmldzxUubHG3kuAOXDKOgqAWsvaAi2e0g1zp0Wo3HPSDp1D2sf16sbJGJ/2iPV32etvE+4XgyLp
4vSuQjUGPnroLn3fIkCXROwWy5TbvqMCrD0V63jU7Bqxgy36kZwHPnJiKP7NCzkbXRQBMCMASA7L
TWP3JGSVvUzFm1M2gx/5jNY5EMG+y1yxOyjedBQIc/Lr7fNYL9HMp3HiDg9gin67qUeCJ6AgdTUP
4LEumYtzr0LkMXeejE5xarePs6ywcku4iWrHv5B70wZj+CdsF/pQFdgp1L/J/zQ14YcbXjxtQ27U
T5edRArHiFdpvsuVEEAElxfpxWXnAWBTvXSSQN6ykWtEsSSHJThXxsl6equDzhBEh4UZXMbfksNm
h5PcriiRg5jssMZqqVSin3svtCrxWhuAu55TDJVmvPTr+OKpEBW7AMNYOzCDmK0CCd7MocrGpnW4
DTNTh+cC5YrnHk0L3fyqJryZVHKWTL5n65uj9BS2BBpAG+TaDgMM+dFVGWlIDbm2gpCYCZdx2r09
0udEOLe3gitvdgoBglpBqPQD5XUq2IC/j0BagrapH/Wdw9y0WyzAA9TNgIaCdc+5jpxFW0M2TVGh
qqZou9aLH2+f2p3SH8cyQIq8nE/O9BCy5k45NPOsFhqKlaS6MuJXomEOJKCuw8o+VDvL8Cdls5YX
Z4yvumgM1gq1716qOS5+7b4yI2rxa2lB2GJNEUlu8P559ArJ+qCNWwF2EwUs+INnMICNoLHKreiw
jzR6LZg52XvuxKUGivTDgmjKlnGIlIlvucuX/pic70ydGliPP05fINxFOPifM4EWL+xoTG6z1bTK
3ZOw35ARZMMwDpiMQxO/I9YZnjIm8/5fDf6Ccjv93hmNJSLZzwAbjanFU3qJ3/KRCDUJwOs3Vkhx
Z/C7HOuVMykTgLYOvVyvnoL5kRCKQGooaWYSXMfBr8Iw2mUvLb0YKr1UImSF3KBBGSJTgbyoDsGw
yGoQHgmEq/CNwz2Lbp227T5gYwqWlrj7hq/aPiTxJlUh1TXZknLUyRl09lSE1i/B6nQm/+PRQlh9
j/06gTBNVI2s7tJZnIgQTOP01FJOy1MLI/5d4GS46Qrfpv9F/8VudH2u+untG3PNXeSIJwpjMqNl
RFuKvS8HmjokvRYL0Ulv7+FPRGEj738oGroiaQh+WHdi0Ejoz6a549socCSaLoi3bxsy8eOwS+a4
RlbqD9b6yA3T+iRR7+MF2tKcJNBLsrkjAKs7Pa4eCxPil6jb0Ud4l9TVhgQ/FIk7v8kzu7Tsf236
LL9ahsH1y7AeQMCwl+AI4mXSEL/6Msl1wcz9cMc284s6O+T/cDq6PjlD7aVwHhRFrpNFihDnT74q
TUbbBqQyJaMVOCqlgYOJCBFTBBALAM1JQIVG2FXEgSmSwPE+S3U7yMfy7zEluAfbIpGNoPJNCcwu
WAZ3JCpHnjt/hJP9eLrrLPNbnNUnt0Kt0nUowtCYdmG/eBZCgOB9Wm1hh6I7MwD76FLAL8TmQMcO
c18Edu3kV6+y7hl+/jiLS3N13TbHYhEymAs7Gq+XZ1SBPkRnBHBIh5GOjOIOGcJv/9PtLVc7vWw/
6FoZ24Shcr3FGr4mEoboDT3x1/GORX9KqZzOy6y7qh3uoR7KeILIxvG7SG1S/cTC3qvODy9zNj2m
2acAu8pRQW2WiGmvOo39FMtvoo9WmTSKbHT9z0r0A0ANlj3nrR47z2HZq7qmwktd9fg6rPiGnG4I
uu/deP6tFB5HSkAXsjdoY+RVwOlrQOg+QObCANNr1dzAm40xxTzaG8e+0HpRHOH8ePEyCaBNWIpI
dCcozdz9dzUEoLozMsYr+6jsSFUh5d+tKp40WjZE8VN6EZJlU950HgEme71H4HVScGgZYCXLvDco
NjWKXS39bBldTH0aVFqh8Wz9qKO8lgYHjbtKnII+6VTqipLJFi+JsUI+fG71UyAdS/0dDCslry5a
ZGRp06gyMsGZFIo5cnT/FIx8WnXCfbeilI5Wk5D7R1rIjfYfbcqycU2oG6WE2RcP6aWddqR7bCce
QmZp0yeKkRh+4v3MBDdgWYFFGvjItP6XwTVjQKCDzpVhLTjSAUsrrGJxrgCa9c38Kn+/YTYTwqCg
k/z7jhDrxenbja5s/wu4412So0Q0fOIu0Ik5eKxqnIEG9etsBCz/KlrYS/J1BYBDXws24qQAAk++
ammabKYb8D/Hw3WPvv0adUmijDYKY32I9OLdZdGLbzWXYLrJn/tbtZRk0LPsNxnVWAMcztMv+Rd/
w9NRoITVuIQ7Wnu2cKHE6KS2G/OmrfTN5AzHj/llLATeyRgKXmFkT89qQlsRXxfcxwmwpvl5oVVb
JXfsI71jKCpvRgNILDRPza/r/u/gDJS9dG2DvrFL/lTJmJlz12bO9Ujv0ayNrNxbIhc810v1XO/v
iwnz65zMFOQR4kv4jVWsoHdU5YHcHQEJEAHomm0JD0BcSbqaH56hI8Wg7hQNcZjGR0VplKPUJKhp
jTr+UETh7OMUNSbbZBUxSMCb9uWMCgxi5Mfqa9xog0GwfVMHadSGu/+ACahT8urtZLkjkDPmroAo
wIhVh8Lf7f6IHUJI2ihS8zdJ/DsRT7QqYSER1H6xZ60oO1jMEyrAA5wY+Dq1AlCoqHzwHqtw/228
mjzhZnpWesTXyei4ZtKr3hkIbwDgoNDr6g6pDGNUyrJquKvffSuQhMHc/1y2QLdgPPxgZ2OhUR0B
vo+Z4H03Aa3Md7Ng4nemLa2vzFDeq1UHvPm/XZsDYdOrgKpnZHr9L9EVNzwcoxXvASgU/YYPLiia
mUyAVAduxyqKt1QVuwjd1Kk1E/EA3VtdvEc8kVrkjNxP/kxDpk5SI4zHXD1DRaAixAe1u110TekK
rismlHu+dmFUGX99hKcX5VfYYu8cW+JYQsyl3j6oRh5gSgDASBtK/9pGm3LF1nFW9oOszOfDnnN7
VbbuL9CDr0925Au7uj0ScQNe2NuhwFYvw7tqN6OGQyNyrP2ACRAdkk2izTeS8W+YjkqG48tTNLpE
koSMpvpXxj/D6UwV6Sa2m9wa36U6arpJCckf27Ix8nJc4J9a0eYSzTzcgpyTZxLV7hYgGgXGst6k
IYD6eTu5pW/yS4hdg4T1CBUyLVckB4DJ1n2A/NU/PkJ5/zmLx86Cposhd83DYHceHlZywgWSChme
iZYs2Nz8AcHsC5cU3yLh2bt0KRnw3114ExGtj9ekQSb17OZpTudqJFGjcfVkRfcWpZbbW9Y6Vivd
sCcAU+Za2pA+xV3Aw07yDcKEVErNKuxJhB+FNZfsvxDESCQM3w2VKSWtP+fsO9+Tkt4H4jcwEmPg
w5nKULC3QKTDSlSUh1qt6RmOPXP+ykx+fTcrX2T3+GPW6cskYojHQ7F5fcYCw15FIW/mpIYJGUhj
B1qG3yJnArbg4jApDBHZTuR6E5esvtaYr5dzSfGfSeDV1MZ4TBq810iChGp5vbpsIB2EZUwVm7La
muGpdNHPO0xPpollIFOFdzIqPCzftT9bF98FyHCI7F5Gx2vMpjD1h7Y1XIES289ff/5CyTw1Snjs
W0TkStlmEAMZnHSRt9Ld3x6VxzKoPjz33lLgBPfk2so7j+pUJCFA/SAjDN6OWnhTnGO+yS+z3Voe
hinOzywn8YsP5R54FbLLY3fxH4hjzLyPO+jUV8KZJIS2xLnMDI8MEzbkPqFsa3qT+ICrU9FMzwzA
P9MDuPH/xJMEDBQrg3gjEdqZhKh5r3Bd1MUirPzloNsgf71pRB1ZNsO5ZCqtQd8DppfDs5q4iERv
wisoyCgRpH7H23P6LgZryQcHCX2Vr2GaQFtgEeyoQvsoku7/KTVSf2R+5/jyyhKXV8NGZyZZ5u/v
q7HRr9TLLoOwvBAcAFglkfGd06eCI5EPlMAghAZ5LJEs2Q3FO95Kl9n8u7qS0JyjFQRa0ng+nwSi
zQyDF7l4tpoawAQ2XisFsWRVnyzYxGipdppGJaeoT6xyepd2Nmjpfcws5gzmocRnFLQqdgwkoFMv
hDU/9S+WjByPMLvyJDTdFg9u8tOejE04TtoGo4poZNCJEF0gTwRjipnPSLKC/A/saIo//Ps0//eV
kqQhDW3vEq7CFYSY2LhuOKrp7N+2HX/arRUqtz4jU5Mlk+vQL3FPzz0/VgMjShNNb7APEwfHjqPC
xI7OfuDk/2G8vfQrU+ykVwGvBQ+rluzDAs9C8G57LWHWXgVyWjNm32sfCPfCJjsyAztDhvgKeP90
svduCIHO+xFLjVg+hZjjzMJBBoBniMVqMv5qgDPdF/weRT1kNSCyeVFdnrh0fi16AmK/vt6OwqlH
JgBHJ6Iy93xcWAgmBV7Rk3Y4u+4vVugTc2npNyvN+n6NAcpLsQY0/ECOAxaBbFdfOgKTmBaI3Wky
lFKDUxFK5kSDUh2KRV5juZOuvayvR32KboMjrnhffJaEEPXgIOW5tN308yVWTFOcPsi1wTL9cLSs
UQoy/vTaYYiEdFcDzoaYxSlHYnwEuWMbnLX2OC2FZO3uLRmkd5sj3XLEUmQkfPS3NbKeMMm6yRIQ
bdGUNNB4oMUF1duy3L/IM2mC9EzgubFx1owggin3eu2ORF9SbOfz4rxdVTRgAlwqVsF2vuZi6PlI
2aVqFvYayX4GvvodOIr2j+KN+jlwSiZz4REXiiqBMtWvsjb+xwxhR8hoZYqi9Fj5GxEF77ejV4TR
7YvGGJFoWYBs3Tr/HUUzlXnLmue1Si7UpiRNOuuobJnzcWp2WiaZ8eXsF6pexVet77InuGdeQ90g
5Co1WzaRaqILDoPmH0KbAAPoPmKM/wRJ6qka6zg+atjtDTxdBDXC5qSxlZVFlY672UjnQp8w6umF
zoZ+bf2FxbboAPVcAndHCqaneSK7jKXbbYRK/QkIbSIdIdHI5Z7/LGaHUUiUOxyyL4FODCby4UIM
1jEIDYWipaCzina7SvMJKUdEb2FiT5UO18teMhxzxAjqsBHBNi6pKhLpSGXqhwK68AhlDBkj9frC
9zrEeYd1zR0c1pnOFAIA7Je0h3QmSjtcio5zgqM69X6ubLJoL3sQwGp1GXFAOPPzTwDLDnLN/gcv
VoxbrvpYAODd5SuoXXqLpkxYklEv+zFHfc1S+c7+RxGbxkxDvgbAgKGqCPIQJkfxYi0JNZkld8Gf
vOAvlQcdug7FQ34aPA+v/3PIR+6Fm1Ab5HWekfXLFP86WX+c6zSgWRlYRnUJ41Rh71FMDfOPoyS0
BbOf8nV+Bms55NbBp92HIKiZ9ssc2fnOsgK64af86Iy9utwpU75rUv9GKeTwDCj0NbAadPUwXG9H
IyytIPB59YXzHHKSxPSwA0CZF3LNd2Zi57JacT2ReEEEoWziHqFfPKaD29RxsAFche+dSz6Zv2qH
vSKgbZgPu3sN2WTD+yJd569Yr0OyF5eT/hiQW+Zsx3pzM5EaB44ueODv187/kofcsv4rf1qFAKfQ
2mSBcP2Yn6fmf0r3yYeUHT9GIN+UscHY39uOUt0yl4+BD79NsP+2hTrRQSflkFSqEEv+/O1IY3gL
0ESI+hGTqCbYt5ZGQ6uEmxWhioYGTw85zIexQk9m2EIYl0mFzeww2QG2tuo3LmWCmj/IbpL+aTIh
fAaZXiUJ1H4YEEBkuRGVssrjM6e5M+RzoTMJ9kttWpnWG013wO4UGdjdyJrjp5ln2ug9OnSos3eU
xO5X5MlkDU97nBAJYe+EuNx/+GlIQTsw2CfY2en1FiQUdcHUncK0KzGEA5Mv/DmpSWkuZJx06RwQ
biESI/CP7hamilr5b3NMzoYuWFy/d+vcMSR5Cofn4+53khOtrGUSW+SueGR7AOXKcVhj3sT5jxz/
E3QzMs6hZw+9xsYrKxiyvPoQxOYZRzimlENeF6BuVI0iz/QfNYTtLo7sX9LiMlPdRNar3cx1ewDV
uACXgOXCS/Oi+kMnd0y22hOmZ1pso/EVxkpSUty+lMmPy84ZyN8RW83nkVlybXetF2UsmFrNrk2c
83c/2VT+3I6geePnmPHS0zTvm3+fCyPHiXioiJqGoBwMiIp35aYeQgjBKUPYj/zlRhw6lwxbXPch
XHAzGBMpGWns3G9tO1i0+3pO8J8OMfbGqQbGEBM0Bcnd8tfa4XBT+/8lmXn4RnGPpwPD67gA/EuO
N1KUh5EYEMQn1Gp3mo8fwgEDRwjPeOHVerloM5zoG/NIkjaXaRWLLrZX8DVzikIe9mQjDmW5DpYa
04mA0yW2AJra1gy6Ja0lLmL2YV3HDaw8KUpTPR/BygW5fVdC5uCBqLCuXdXAKEMssz51NODnRmne
yQAqFv4xYDe34Ql4cMgRKBjDtismzdmxjb2zaro5JOBG4WiboVe62JCGZPheuasf3vlNvZ2/S3o0
hFa3t2A6u8SQ+4dumnKHgC/01UNM9dKRndfEpjWTKp9GTQ1J3JU1qwyOmuRBLphOs2IuajRnoMjx
/BnKhynE0obvB/WNu5G/Rbry4626pfJ8SS/bYP/ChF+8pUKSFyp7ElzEPlt4z6UgQrbuBxpWkYwA
TYcWm0DKsHOJYwERRalXCGNZIcfAqp6Hb6urTJ73KLnaVenlXITAh9rJ31+y19KJB5L+3lHosNZr
+9O+RRJRab/dHGiYbbBkgqfb6RKLtbqZ7TBdH2gmF6NrbbAjoKm/zW56HYM/qCv3wK3RugUkYQzu
bfM7nYglTwgsHB6eePxNENzG4YM88z1wD8KhW4Nay3cMxmuDRaR5NWcbMDRSl87qmfPCjIWDyDYo
BkoXxeGcmHYWjbTmKvfLLzDtrgchHLPFGmBFkt8UiYiVAqojpsRuefgOl2Ndv3Jk77KTEBSF0/VB
2z2hA1O9Lf7OXmpHjPQc8+tAnVzMGeRln66BRBDOvZL3pCgKVd3bsqgH6xQ1uwBisOAzl81nQALM
9In9z+tqUiLdvA72/IxksVtKW/QH3RT19qRMHeyqJHuQagIvKlU1/plbkiTvRjsiso4IywmmqVjX
AvFGQnPGE877LBu3eLytSJ0Xi6nlp5xJGUAB2TDckdjS1cxPqR8yhv1XKOce27OwZGD72mfSkidR
cSC1OmxoOetz3xOdWg3dmNJIs/959AM3f/INkV1lYXsfm4Em8OfFJLdfGvk5cQA/hKfUReLI7tbr
AN0/KKB4P7lxidKdEN2EMfIgUkmDQmVK/WGWYUqohiulATt6JymfrjqNQiRPbv93lpPu6wZhXpvu
rrEmId+kHxUGmcbjgz+8A9whRp3kQXT6g944Fx54VLIsi+s3+c4zzM9xUkKWHLZXngCd+wXHRlW2
ndXFN8w6myc3YdvLzASE0AboQTw2uuXSQrr7ZTjd+rv8yDBdE/pDJWbB3gd9X7LkihxTaLykIBG8
Tc0Az41/hjUVMpPDn8grrgnqJHyH+UV8l1gcGpR+P9B/O9M1dvE+leEOx7bRX7iFuhQAor8FYQNc
smQUZ0PhIZelkCe78NVVVNaqhiXmnuQ6LYKKkOVG7UNzQc38yiWwo9asYnsXejpmhrlIYwdA61po
3FVtxFrtXQ4Pf7LWFj3c4iHQ7v1yjuYU5BflGyNO9nrvF3kbK+8XqevIBMfpmVObFmh5LXh9UMDD
aNHmUBX/KDIZdQLMfXIfxhVPLL2YMc71xV/VbpIwCwiBgcxK9wQA2bOdWMmIEBlFgfhscvAXwqyl
9M9YPXIgul2B85ALfpmdayQVGbj7RP+IShl5jHvYgCVFDRw/MZFuAq8dRBv4/w8Et4ykh+VxdQaL
lHsxydqB1xba0XwCkc1iMklL0kn7yni4xfyr/BSAEmyaRh392euv3oNRAgxhyYsaFUxK9e30tu0+
jpLTOr3Q618NnGhOfCiYbTwykWprY682jX11pVjyMkmZGIG+rBGFROOYMbJ4HC9ndxDfsnoMNzZD
Uty573VhAHVYtGIuEwxIvD32WgBFVSripPQ0DgH6y7m9JXPIw5UU9fsKnQP4DxelLWEJv6MTefYG
eaq7eGwUnQrSYoFH2ZLarS9PkkXsFOyuX+PuvEh7VLwWVC/cw7yFQk0/JILJ2WSskD+5ib+zJADr
vaqqZHAreNdTeLsv8qRdFzsEdPWtffBSFTaCyZUilurXX5Ll6oKcYwWalFgFhvSxDpQQxbsAJccK
sTh+nqVzBftPVwkjoVZBuD2Bs6b5RKnIYD5KkHjRv0ZD9TR92+kEQ/AzKaRl7aWb5Ucb8MBISvMS
mIlPYz/AjENVU2AEw/bc7QQNc9f13FrHwNpBSp8r8c0m/cdcUDygpMHjKN2J7blf3D34XyYd0dVB
wyxPPqFlH4Mv6DYdI4YKu8QrTIs8m+AlHDsHfF1XbPWmt1kAaV7DB4zliDTo79ob6uAUto6xoJMN
XZ7Kp9v768je1Lw09UjpQHhxFKARfmRLoHMK9Pl8uh7fiiyOREsXr8R4CiTCABk9pLFS6jLq+/zW
+vuniCvqNvreoWb8DpBXbXifFwXsRiA7fJB9h8m6CotgRWplnjYqxJzsEvAXsfONvOxG0FLDNEuV
NLwuCiYZ6sukv+0+RknPpSYdjh9Ag8yiIKNI1ExTuqNTGBJvVgtT8IdCtsirMxxu1ePp9ZWRGfE9
6N9+qiUP6onE6oMLURLOqxcwsyE2ELUlhevR4w0aJQbnLt0pt34tFks18WJjo1Q9PpNf5FluIh4F
EbLXyFl0GAyMjpI1Eh8l3LmEzu+1/cg/m+55mA3s8VIBzw3MsCB8NLUZ2/wWjsWuBLti7Bi8KJJA
ES7oRMwfuZ8CTNI0U+fjGT/PMUtF+RjSOtigOIrU2gXO+ynAFN7GOPG9KIz+LrlJDXwsFF3sNBv5
Pzxx/PZGyQmTzNHq5mVIjKU40/Jt836Ky5ZOWWdvOPrqnywbskzSiDmRmEtk7MrfkQdcJS3EiF1X
bzZ2zdcgy3eEaezASJ1Yj+Fs7hxb8bxt6jFwNINk5HpSyGBLuKzAUQESDoQdEuodOtIlxUKfYi7D
W3Cyp1JY3XrTde90MR9McrMfSyuCe5MW3Dq5E2YNsfQjv/0W/3mURSKfJu37iflkxkxZYaM2EHWB
UEPfleNRzxwlcw/zGS8NgNFQXDOXuTEVxivVmUcxbpyayDbKpkY9E0xdCbsTTIseDWLz1kZlWl4C
GigptZARuRX3bKhjzJ5xyfTayr+sMyGmmFjE6UsTDbfAczrNrZe6BahCwfxxHtfcy8qt7b3PlqnM
Pwz1lgQOcQAnYC686KxaItm1kna0c2n+jw0UErO2YSLg/RNTHitlPY3t+EfQhZoAV1/hzB8FFC3F
5Q74ydXvXaw8pl/ZDkLDW9OrvsRSLrDDfh3cme4rf+nXRZnHa1ZZC9/yuqVH9qDhZ1Xsgyu3s9SC
Xn27nLRbO/v5A8ZALfNuVysBqP8UGGC739UrSCxfsUJbpxtoVhV9RyRmuZbjZ8lbQI0mX3VdalKk
JWllC8Af+lQ8kkJyn+scsIrBWuPKKIzExcXdM73fHMr+wpDVbwEPEQjVbm1dqeuDoB+Msrqa8lnl
Vn/AIpjY4eQwO7jRQ8tDieCFHwEdU4GyGe0MgX+fysVGMuEsKAp2xEyvZKicyGmPTMLZAmohA3le
2Uk61gYMVDLhhnOd1JjWWNZ5r7RiHvcO13a2X8DZNIary24Jo5aFa+c2ilVE6Spjth+wrC7bynmF
FtkA9gwlkGGI96mOFyXxE9mdwW5cXuWY9PqvtTXz/m7vz/60Nph6ZetpgOlrGp4f1wZ8rtmeY/Oa
tfnqiGJHF9IkaMKTD7EkDSZB8gzrYKRod5wvphLVkq9ATRJLei/LrlMNHSIFvG5UwaAqAQY8NRNM
97fYt7+otMZPX0zmtnIsFMJtHsJKOi49V+TEe8sGjyVDZqDSDIUTv+Fpw8Fehh0ucjfAymIleeFB
lPjHvRv/URX9G9rcvCj2gM85HdadFPcn4RoQ4vQzCiiNTFMj66n11arxzCycK20q/SZA5Yy5z3e9
hbZHkZFlBVsiTWC3VPPeIQU83/yduZT3Qd2fy6osR4FqN7AtsnzBbPjG9AG5oxqmUpno1mRGvJaf
h/E9t2GPQpEKmuKlMdn25H2cUF0iomd+r8us28yeC8hJG27xTdOpCMFsw3wG4Gde7Q2rROfsvgdH
kQjSDh5IkA+VZW1lq5lOrhWoCmyr3Ke3iWuDhk1fVRpi2cV5BoZOWwFBeGR2VS5VRKR11zOZfpnH
1+EXgoih3KUjEj1l/qLWgQa/gkKEGNLGB2/glKEvvGhYbamidyRRy5tZcnlENlIfbT0TpLvvDD3x
Q7a3rxNqJH1WMXm9TaNN7kUhWZDvM1l9Ib5/2xlELBrzLHod9PucSrltsih53O13LQkq+MUyHQ/O
1Ng/fvRb8febG1ObH9dIdFDa9IWOrAm60xzG96mQuSSnMhLtzhTL7iMWOt0C2ozNwHGOFJ0usVBX
27zLjnQ4bEnMBoodwg1iBknVGRF2FE6dbBtLzyM1FQrEX7MqHTc9ojTCzUUhyw5ylBvBcdVoOYma
XjvFrKt5D85WkgOzMcVhyMDLwQ5mPkfGvDBrFBAF5h3UDhyO+gjmX3F3jPg0a7uAkSLeQ+xipZkT
/TTJ6nC1/rKfeADyTP5J3tpvAZgS76nZ3wXM+Rbm4TscLdrla/odAdXII4Vv6bufMMVP9qjpwShk
/gCW2FYZSCeghmudOGvBGEgkKYymDZUhQJXp8DzmE33L4bKHL6r/kVL4EaPk9Q9z1s74E06fgKS0
3XYQbztFFCKr/2HM3Ml8M7q6gnwKvPfRcdDql9xNOik2xQPCjETesgDfwilikwmRneGrl3bC4ZAN
DY2D7ADlbVZ3H1nZAcfFrTfGEOYJ1mx/yuNug/0Jt9Qo2HjLobUzIGkk0iuZLltxt3HKr4u3zwQo
L+OPgahc2SMtQCFpNRRWR1hrt0KLFjKaNsI+XvWrNcVdR1mrnkBTCGDuq2a5n/ihogKmIgfxNKIW
n39pldKInN0YQOfO3Bwo+uu8sxSjXtRG0mdUaKwkDDhz/iaVQ5Cg1SPvngAnByuWL19aNo2w+5D/
fevwuy1ArbwdboAGzMjzIpYGNvyJv04atDYi75XoXs1qSn+/E+WBoLd8XUUiYS4Xvb2pHxrcCr8+
93WI/n/tWIHFeUHS+oU8s0+n+d/1ndSJiYSS3EDTjyd3LiTEz50WtU/uPg01BhzgCyRJsgX5k7rB
P1pOrt9AFeHq7DeqXOXTitcYQYnXUsEp1eplqLtLjTWRfaMZfd3TqpgzszyBgRASZh+ToDC91JBp
rx5x5Xl04B6NCyZOWiRkIhGCPmDRfliqjA2lmBP2YC794S8jXImGVz/BuJsQo1d/73ykfJ1QUBpT
eMLMMe52KXCcRzWD7XwMGCKSWf55+YVCn5pzkMDnJQo96iGsKDXQNWcu9w+ksQyM8+XvIEaUWxNL
V0JzQSBT+Gc/0pu8do9u8D+joDJATLtJP73Gyx2z+kF9oRB9siO/aPFouWZN1VMJsa88FbT727Qz
6R3HhujujyZ/soA25lv+UhSgnMN3bUqitmmoBnJ6e0r5CvwuA+4TiftnVZfp78OMheUNSj8l9vPm
YjSHCCzcHD1Oc5lMM+B5jyyyWEDllvUGTCJe/Ue6gJwya6BeimjIL1OfQTA59e7tuFZtfWmxN62P
GqM5SDE9lUmT7DHdIRhmQPU0fjbyKC6mdMD9Wy40IUrf5x8R1RyzvypFu2laRdBSX6H2ppAuEfz8
NZiL8/+P7qWuRbu40o8+t9mzObNUP1ZitIRlmZl6zhzD9p6c8apxDpUWXcSxILUSvPohbWZyn//j
7nHNmZSFAIgv6JUcvtnsmfWz2xM2KJunjdG9JSLGrrhSqYYUaP3hkHd+IzHlQdJq8YHEa13Mopv5
t8wyq1LzNM7iN+2woddG8CIO3GlZSp2gmONreSZ1kB3Az1e0qWVixpf1iP8Q8ZkZI5pl5+vMDx4R
pEZxxHviYufKpYqFD6GqjgRxOjKJHuWUV/W50mz5GBwUIBPsaYoaItgvPEQcOKq6/S9TnBXQTVrU
KRZLENrIq/SbNc81t/CxH94FU3q3mL/Ye3dM7r1tAaZPazepCVBUID8FlqVAW7KFJfYsiRZGaNZs
O1MTV5T0vZIWC9uLTZgWxqxgh/A5mhBuNXFjA4TsttizlTbpDq0/hfo23s0oCmL+MA1VglJnBNFe
rLdm54q2IveG5Wa2bfjFm4Z7Ue5mDzSnKwlfr53nWvEAgaRpY7u4v7hN70uikmsLszNvsL8ZdDj5
IpIELSUqQEdQS1qm2XbzFobElljrQBToYJ/jX7BgZrSpk8uX+M8fHjUBJZldPqygy9Y+L1U+xl24
AreVwewhMBWZY/KFO/gHtHtL7sTB5H6AvwbDcGVrW+ElMZtlUSRxrBUxcxXDdSrl+osorW2BKN6h
Zx7+FGqYYjtUXefgGZTJ5swqr30R2DIjcep8vCOAwF5/JDbQZvSXdmfZPC+GZ39DbxSiVQ+BOxFC
gYHrFGSbWTSnIEWLA4SPxD31F43IgDOYCB21nFAMVaAzpbqVu+3hbhxk2SbBL1VuOQzxx8bkCjHr
Sdf3OAOm4CSP3gOhG51uFFR5L8N1CwYTgqAY2DrMWUE6FcJnrUAqkjLjNIUruLj+O4mTrj64Qj/g
U7b/A1sgfyiiT0rDurULa6gzmfQiq/aa5DnvL9UQrhJ1ZBBRDQ5HIMfGhAp5vXZMtWaaWXVKts9j
CvV6t4GV51eypnFhiWRJunwsn+lEaocIq/X2z2rB2G6wdHKpgTzouJN3z222NRnRo3zEgxoTCYOK
3Db239aeqCHikGV7Q8oLdpdKJtxxIzUCudgk3NT+GbXJbOnx3Ay0AXphpkUAgc/rOUZLXnZzDipM
7KVs7yEOXlxkvkFgKwEanWCUPUgYc8cseKjN4CpP9eTKmxOzdNyKIkt4hjxkbQoYSP/UNkOGl56M
YUqxoQWQlanZeW1QjRGc+oJEMd7M4tPLFWa6m0MjRyljEFWfU9D59vEjQzr3B7IBZFreefrdYlWo
YUVPT6gWH48opcRBVZG6bemmFpnU7gKNSNgmXYmou+Newk9RhlrcsW4At7hkbgOWqxzQD2vQbOPi
Aq7Q728KCYRnTi9olsQb+sDqdvLNz+r2/YTAhxWs2M9clFH+uEy45ZsL/7RChfXPZNuYRDr3QddS
kmOuchoywxlS2HfNOhpZIZEAznNSfnYU7tynUWPTvl/ShXemO0UiNlB9unAhrjLf+d+dpniVfo5z
1URyxKLdl4jR6OX+6qOiI2B4UHfvAzphPcTOrPQFLeUwismb9vIIfvEgrLwoWDNeOGyLfUhLWQ9B
LllpwKYC0eeCoAj6CqoHNZ44cbuOP/8Uh0T7vC0BrKITQZsTUmwxiNBCg+lJ+RcH8lt/v2iyTH1x
7smaAjdDLirK+JhkiGil1PTCot3bYadtGBW/4uS3/LhPjB6WiA3yf/C/wrgvTI1FcaLCpBmgIPNk
ADGMdq4VEtvXqCr+910DxE6LPOuW1RkYY3jsmumowT8taMcKZ5sWN0nyGGjHDydBKlAtAErC6nEn
eme9Ko3t4ORd1WwjYrWelxf233HpGqmuQjWacE39Uper0s2cR5kZuIGfXQd8/GSFjxjsa0cBOiOB
ouklnoC+Lt9x5PsZqlWOereaw9RLnoTLBHy02GBCoMs57AYETp6HhBCs50l6WyZBlPihY3Za32rE
IsO9hb2JkQ7YNtUp177TXrPblEzi5ahg6pGKR9aWpEDe1Vumaf/EHyAgUzsxLAdELPcmUf/In2My
vyBsJR+5tDxsIDW0/MG/NoOGMB88U1w89N5SmLi4JeMMtuwnPoMEGY5Yfo8eyRLtprvpqZ2vzTek
Gm2RPB1XkfEl759PTysq08MCp6QPgsoYC8mndgwdRBH3a40/qXGsmTITG1kxKBgZMUqf58nM7J+P
5LNnBv63B+SaGdKzjxqyAVhaELTh8nO/pSSpuwAsSCBByfpjo9yX2fPaNlquf09KAUikdi5hzZcw
3lp7dPsxsI6aJ7I3+jQRhCsHITqH9SLKseqC/EkFcthxdRCQ1AAtxYRu5thZmMq8yREyh4bKnQgr
zge7KhhyHLNxyOBAzoQgO0Svc6wnOCiVWgETY5S/e92qrYdnkHPcVBulogPCWuFRL85GUy4p04zL
xMMeyvosAOUG+uGPVEasUqsnU/ot3znYM89v9aRWZSA0hepwgWAYhWxhmoxiliHiDamO8QaQAKpm
NhIYJa/8VVxSZnSVNbGnXsX2KUhLuxSfv+hDQrAHAMW8/uJW4H8Ij/CPIRDcRTFc+IdhHzgYBfOc
UqQ1VqQ7CvFt3e96HD2KgJffEXXRzcpa4rQqJ909IZzGgktic7XDhXxRfJlBsq8bzmMR9K7stNVi
ERqb2aijFksCn5AUAEuEWG4Xcq1XQ26+Hgkm7KqAay/96P3yC36wyqgY7SvY+enDrVJDu0Q1VEPI
sjSk41md+AJJmVqyKX7VnPdXoggpaaqtGTC9LVQ7ZIIqZXbAHjqMnJmiTc5+c4BehQsXMwuI1fdT
8PglU245JoALxV0U63iPHh13f7XzS3ubvoMySiN9rK4W6HSduIK8E0XL4kYfzjo5OBSeYqQj6bNM
4ay8ykMEN2faVsK487a2qAp9LQOXMyrh2NAS+6VsL4KzefWddy+H9tjcxqX2qpUEOgW6ONC3coy2
m3EmF62Y3FEXeSqSr8tfatyZWWvx3vCL18q0EhsU8RQ3SwDG7ycOAriCJDBKR6LEE1Str62RHrlQ
Ndhq3ULPNO+/8HxzS6XtYH84XdNqZ9jjOcTyKlm7EbiQRxj3U/AgAXK8jQS8wOVj1DqJl2ryLafw
G1YydeL29CYEclq+Nu3wbvWwWif/O2IlceUASXwTBk2F9z808gH47O/2v8JAWjwgwhnUyeMskz/j
KWgR7UETDWqKmmNKoo+1EIESK3sJwi8/Pd70vGT2p8LwpDJH+011fIflBfGieCRBtlLs3C+IpxHb
l+XqV285GKzHEzm8SOFqbIkxmqirK+N0R48yLc4ty8BbNabU24H4A9+4P9KiGtxp+UDdqI93cYAK
W68ESW1824UYVz03wByE/HWK/DsSywJ540NEriFo6cVEgaBmKPPUx1J92boFMtejAlbuaWh+ojyG
3yQ3DVWA0GB9p/Vo5bXZeVhODri6/ck330gU0uBa69tLuA3ZEhfcWgyuNcFCGuW3M5BG4xroyyHg
1GtYiEIcbGd2nxW/J3KElv72u73czgExq56Qw3eUb9XQzMQca04FPjaC1LbGqDWq5ZdO9z/NYY5z
vw7skIctB66XHTFQ1XRMAipw3+j6y/PKOEH/RGewKA2wDWp1qqagliBMWJzUpi2l9AIVaY4jSb9z
RHpZiWjB4/IRNskhSCUEMbJ2G19aIk4w9Jk3EBzDLgpJxErinajIxx5ib7P5JKmWD5kC4SOUR75S
pIo26uxIheFw0DEnutreVVmrJ/V+do0AUoE9htLkzpdAigA6+rzC3c74AlosgjRPY0QsUEfSb4ez
6VztiJBjg4qikYdUxt37KEcLJPrCQGsWGv9qXIAGF40JIUqcglrm06q0Ux9JvZWMNepHFL3qpspB
FdjfMySy39ToYmlidpGuIAzQE2wJuciUbMmR65UdWeYn17tqW/a1+/FCyzZsRwIajCJL9XKLi0E/
FIivNTZ3v4ot60VVnlRpu35IAsCpyiYoSjh3AtdJu8cGO9L8fp2WideI5+mP2lO9Wnj3NEXfEga5
mcITqhD2rkdJm0H5Aa1limzNOqrM8KoOVOZtYHpaCSh6BHvhx0JVdxwqywUYlxCgz/C80OePB9Ap
A6GVGa6ZXurKmNIb9+BZX4QP+HnFKWTqDJ8jFzSkjPIbiD4YG37ycXyfqrCsjrs/I02dQfYRMQKc
dfMeUWP/G24v59eirV5mXTZJYWknR1w7zDhjoVKGuvYznkuCjQ9jDhp8cVl0If3IHOcSgvMKGSdD
lTb+HtrBx7NlXtGGy5bAlPvemW2yvdjhfY4D0P3rLHr1Fm3YDt8AQ8MEvAA+FbzYH3z0379COZ95
y3kuMUARM9Szji1wK9jTzsBQG9DPhFvXMXl4NC49TyoxY3Wq7GcM46ADzbkdVa/zWZTPBnG5nzNS
S+emXtlCre2Yugyd0R6AKnLwZW9pB8Lqa/scuQIOl4XFG14/id21tP1IJWOlbt0I7ikpQwgxKgwl
ufol32YGI88hk5j0I+LOBI+ceHYNHwEY54Bien/2Hr2S3vIn9aI5LrBIUST/DPdOyAAwf9mWFh9E
/KA8Apl/bEktSg5R2GnTsieU0GY7xnAemfRPmO210aMQjTXRZZmzq0f60lSXYDvUMjBcNMuAgA4q
mQQLUOoyAGDqmd6wk0//ikJhhcXWAmyYb6SKUYMhdsKAAs8IdDMBpQKtAcSWv1JYEq3psXwsihht
3NPIcDIw1KCPU2usBHfIKxDlx/voESQBF8fop5TQKBmNEJG+JLi6lzbXswy3OzgokU9VQtWIWAtA
Bbdcxmgaj7li/VNgNje/YlZ+vAYV76y+09EVSrzBx5qX5MXn01rVjIcmDrHUQltzwzhwrZgxKUFY
MxdE2kFsw7Z/Q4vp0RwJiVsuOr6d1DuG6elTESxq6vY7o6F+8TjK80qllohQntkgVI3C2Leml+Ps
InsYIn9vJxI0QLBM6b9xXhtF5enIZxIuYW2DQ8+EDzDWXWBTC15uT21XXYwsZEZCbWLrXrH29ROX
TUj1EhyIwPJCzIIleaA8j4S8pSWhkdIf8MUUhn+p+Uctyr5I6ERWo7ZGE7zkOfHeVSJP5NJSxGYV
EwNG6LHZw0oV95J5m+8R8gCzTWOXouoeHWp859LFlO9swRbBdjkM/dxIzmPRfjzxiGeOwmv36H/q
WOQcJeb7BthZMkTmhB4SzoMCu6e6icj6BSoDg0Ri5u50rtEbP1iicMZ0imuDJ/hEnM+m+pCqoC7s
+PAe1ktbCP+ET3R8dxkINsZnxTrXCWeRb63GXK+qtYngkarHvukwDRSbv1ogNfl9u3apzrszF3AP
Lk7WQUaUV11cOy3EdrOodTdMmNXPkGgCSARVY41VHRbyN4Ofu/4BJbESDQd/Owzq7UXCV0d2EqtE
S076/3QaBFM31xTPNKT2AphK3OkaTUu8TtUIsO+nkI86t0yWHLYmV4uSGaF82FyoU4HFH4aeF2oG
E3cnd/Dz8wJ+ydNVRvSMEQP/y5ALeN9zPWdLH3JQs6/XCcKeQDUr6YUrFjHZKZQB3p7ZsD1VtHgz
dt3JoIqEnGvAxhBdPrvV7EjMWwHiffgV5RhpLkf6f3Zc4i0LfpzYROReGOfqNWCfSYocvjGzS7td
Anu860fBljnzBC8TRkfQQXB6bEISCw4DvRYmT9fGWwjqPGycojBa7ba8ghxEnsceSfrMq9qQBFCO
QjDGuy8F/23X6mKywup/k7A4Yxtqt66jI8zPala9r2g/lRTHkNX5b4YppkY7U5rK9YTavUmJ/rit
ZhzD/P/gkIgYKBr+uz41LGXe/Qdoc4eZbkPcKNyY9UqP/MCDWncEqIynSN+sAyKZwlAp+5P9SYB0
FwqgxEo0rVxFdJiNGw3xeJtd7Rmw8ywO++cPiCy17ltrJUOuIMGvL/o8TcXXC7Fousmy7bB1iEhO
OFTIW1Lg9KrfovBXGszXrlBxt3Z7/HHDpeywIDw8Pf6xP3DX3vQfVwHe7nMvJ7CpE2VZdQt7PEfq
uls+xN7us5qSM4JX4JA68vB2tg4xq0k4o9Y0k8zqUF0TKeGN9cqVodpgsEUDR1VyQlR5xlbk95eZ
snwUo8nopBoR0Cw9swwFmYB8EMIJ+CRA8PZUkD5dR+8aUjRK5qyx/g71vcReJo15RCpFywHJpuXK
9zu4CCDXD8B6njEdyopF35owFZ4483z4jmnTyoTypVw+aCp9T1R0Jo8D1tXq8+YFFJIuQsXFGD5P
BrUg9723w1X5boccNMOfFr2uuxFIonb49Y3Ob48a57xG7tfDfTITIQiymf0FWoHkeVhYgtD1/fAZ
rbZzrz0tjZzIAhVEja8Ntp7ZnnWVXT123hUkNImzRW540dKAd2cNAbxoEGKrQCVIhazQwWQ0LEEu
kM1cQnjmmCQqqEbbz9w9r7NmUsTdPPYj+dvSparO9DtWryd/9VxYT7fL5xvT8XHfvJmCQrntarZt
v+2aK+htAOEvo/aOteRviQCNfVEoCwwSdw/HuJhAaGPL1hIpXi4hN+oNQUd2RcCjfVHFY1DfoRT0
ptyh62ZZi25I4AA1HL4of7O6cVDVFm7+O8yWqkIHqkbyxuq+MQeVrjeE0EYf1l5HVBNvv63LSFNs
RxIadVZ9zJkUGhFT5I+7NY7DvTK80Z3J3SMqyzO/zLkBnkZxTWOUaBimg+69kyjrl5XtdWz8RWAT
Q/tZOFygyeoORef3nGjI9hFGPEiAuw4J7rVHIc4ylxParulsPSGt/l7Em44QwHiEJkUhrHEQ0EKM
HF1DdKbzPc2Jd1WQCwnKYSm39oL4GF9bOMf7Sf446EvlNnD5U0zJCKlE8Sq5rLgOWbq7e+pejD7a
2UHk2fxnsKXWETm0ird7Yy1IIZm8YXmw3KDo4MHpVR7re4vB6efFiR2VBGG91ibukxHYzB1cVnp3
DXuvNtE6NqBXUSEWkIKM6vrhqFRegV7pNL4jGpV2NFHQb1RWYjO2Y9Vypi5Z4DZuHEVXV6XgxQvU
DyyiPW2DhW42i/d9upTzTLFQcIr9PtvOwcy3o9GxwAwOwYnfw0/JKv9pAF2TnKi+LpaZuhIh5ptp
5LSTujnElukafmOIM4CQR6AGRyr9OnxsZCFpNzS5JQLhxlNsHHSxyrbdDbWTfx2kt8gfEVlUo+ru
d/YJ8tWhZpKqfdPbMRt8psBjYjxj0HctviZOrP+X254CnayuEfNj2FRc4LFCkLxLSaCbLY2REdhR
H2NLZwPpBL9q7UmNMrkgLb7GylW45hP2JAyj7SC1DFs7gYZ1lmxqLPLaClrzqsz3tQ9t9W5lo+5I
GX7mW0E2mEmhOHTSI/yyWxk0TkAWQ2+NINrRtXAvh+3lcB1+alxeiGW8SDy8Kcvu1oy28SJTg//8
ORfljFDBUPgX959BMw+CntCcYTppNcUVS4+cjtxQD3HIS2kCSXIUSk0+gipQF1hU1nyqTugE05kR
WR9cTdSZrDCL6QnLetRnhh7cWiLA4neWkqDziEbf6RdU/S1cVP3azibPLdg7wsWTKDoXFYu2hUnj
fyLXXKtScCBsc2ZsyrAYQZx66W/co6gPiCwNLBC7FCrnO5ckqBz+P3KlxuYeDcf8tS5OeW+iW9n+
Q2TTQvBPB63PFETQB+tCVbpK65Fi5FZqnH7jwqxV0DjroIOKFjCQvLr80aEm7zn9Yx/HkBtLbdt3
szfK2Lunn13i6J4+QSwlrYNnNv9wMGTGvsoVeWOWO2hSRFeS/rGLwvEj0lgmM/rw/yj/3mWAC+8l
31P3JRdEkNG+Yoo9DrOwLqrTFnv08Btp1dBkSOadhk3hjB6EKkilXnwxtpMMEjzHG6YwZgm+uzwe
dIJq5UIfrIzE432S68y/2coEOFWoHVXe5TLKC8ZcRyoH4RFbX2wet3goRDZ1FjRNmnj8kzp6C0k1
rJc8ZJf96KUgJLliOLocdyNVJAxAlkJpeRvxu9xj4uNW7MJvIgDBQtTj6JvRX41QWQFQkLqUrem6
Cil3vekiXxJPDa9eFS9QQg19KfYnfZRsC6IuWKc+BzxP+QChFNUIj6EWN7E1kIIPezqiryXiu0lP
FzcCG2u5rLkq2LlryX2Mi59VxjO5azo5RGYM6t9az7agaZz+nOUdbvADCuhTq+ETykVVDbPWIixi
zwfmNb0DDgOSP+WoanWKCEk9OYGqh4NjuqDvO2Em1M8wWGwGckc+LG7Uvragm6pUGRsccyY9XFbd
ZuQO7sU2b105XrmNmXycTJslLiw94cxedRFJqRmi0F/TskdHBoaQYFEsPN+sq+GohsS9o/GV3XId
ouF+iamW3LySD9VYnArxs40EhIDbV0V/4ONt7Cs3lYKeiik/qvpRGxXRweRmAnjiKruwU3k3sZl1
LsyciXaV2JyqM7O96/KEBIfzxU7+kD/52wGZ7MER48gNfvIrG0jOZZ+GwShrobRahegqmqFt5m/U
NsA3QXz6Ccrprh+SqRjfgUjLsbl7DJzsTVswtxEMoqknV9VHxfurySRWkdtVmUmNTP76UaKiBLek
TQ/6edcN1DWVLW+ymcvmmKSh2CK69Fpo0MvNF8Vwo9vbwRTy66Vgd9KxQ3EMb6kyAENqy3+Kfokx
75/0WdCPfpjVLq+63WKFPEiMRb/eG5Dvi0h+R4VaMgzXBkBh2/OunoNVOqdNyq6edzMp0BdWFivP
x0JcyvE3JwK+rktl2BpL7o+9YDmRmCNfgIthhJpWTuAnOehuWYBPzpR7qt+4uZtDv50lYp2C7VgG
JouqGlTFq0bXG8AIbbANEDLXIUAiFDnEOL2VzpI3g1HRK0UCmkBfTSs9T0b+LZMATxTt00XyC7YY
c19yY5B2dWYzQB0+GS9msDIXGCWire6DTcwkvDtEA4zFVtGNtURQzzqFmPX+W8vJVj9/h9DGegC8
LD7ust328gggRo6H4RmRTJbuId0FfY8CVLLpOhRTPE4Z+X90BHpeNLhGccgUpWfc+UIBTZVz1lcH
V0sAINY+Hxt+bFma93juV3rwNzsECa3j/lODlRXvKvvQW5CZ19jDADl09ACTaXHwfrxt9UkwK5ZZ
UWq+Jxltmky2zJCtoblHfoe7pcZndbn6GZ8RPR2gFGf/1AE85+RbsUPF8m6YbjAjMTScoJ1rHfvt
8l+83aVoH5MJ5T1lqgG26FwVa9N8OawDDaZFH62pMZ0KlIIEK9W4uo8nXjrOiHiu5rYaBs4jq3WJ
Eu4q/vc9yVyGrMzhJ0iiOdVZmu1bAOXQEP9V6gvFOqP7whnhdy9SnHPsDngoJAI6IZEdAd0MWOJf
ZjvlT+tU8ZU9B0l2sdi5EV0Cbw0gAfxZ6HPkSx59aXRyRSLERuyTUJhI12wejhg51JexpNmJFHCN
+Isr7KMJoIqwPOQ5f5hUjYAPkEo/XYVCZXRHIHkR5FOwqrxQRFvXGerdZfuAA8BRUulmqqrB3/jy
UF/DLR7N2K59pvWYSYukvtnFs4/f1eBdcfpEONjKBJJdvqC8E5/s95jNIpOdgv8HDvl0zf700SPY
I+zN4oOVYJkvuzE6kJXsjzKHpsVRxN4ftHPaCa5Yw2bo5uPO5nIg8m0ID4kOck72ywn8Ai+ggEI2
1WBAG1PGRiOyyvwSATZLbc2xYNKC/XqWvj7Vz04wWDQGbiH0C4vQINeDRko33BhYG93s0SFrjdo2
Z3ABepj9DywYF8YNnoOgz8fNf5GkM6a7HF7krxgHJewYZo5o0CKVohK30IRHvHs6KMS/RhWMwM/7
IirSC0W0scDU4rWilHt+z4AqDjcMyzXpztTgv5aEWhLVwOeK49xyM3tvLe0WnpAWGyXtlmV4btBZ
H3hgy2a5zQvktWLge7V+gD9IM3SFtTh/13Dz38RIqFQ+koBwsF7p0zUeMBuRxIFpZO8QwdYPKqoN
5/f63MJwXKyVyGSaITdJeeUSzm8QMpoKs+iyV5macZx6nZoVj/GuOF3vCxisB6mx+6NrF2Hv5VLa
JnT2j2ruRIbZhGg69OPDa8zbSoSz0OkJhH68zh+j8JWkrUCWeLLp1DMypm53QFS7xL1+KIyYicqv
UIkAH4O/AYvm5Cm37p33a6f8LHrBT8tJGazXsEvnTpwQZrq0hen3JMFbFSWlQgJcPsUfKpNiHQ6w
lUDcOO52RoBl4hztOr2Fo0UPGZ+tEmHqgXbQdrBDcPFDH+Gn8VhnbtuiIYI995DqAJZcCetoxMmJ
RoumrSp69tG3tPySVCh2e5M9eZD7HGYMtFD73mSQIk0Lt2a79PUK1S9DBz35kubZ857hJLnkMMvR
UJ3DHclmA/nXHI78atb3f1P3f7T6JG2Y/ZKFtqddwjYTLdb+89/YwIjjR/vE0+iRdb/t9QW6bLQO
6QuuN+ESIQgR5TvVJu6DeS28u5jW6nvwosOm06AHHBHLKLkVNGiceyQLt97iboCev8rrwiTvneC3
1mwI9Rs8dXU1t3/vtNjHFFCxTGXDazk1+zjeodbzGQx7+W5Aceauw4D8T1ADnzA5RQQkWwhTmAMs
ibsxgmiFs99zOhQElq3GMzz88W8yujxd92h/bHFh3JDtHIdnYkITlcU+vVZXG2KMv1SMD8rck/cP
620tFRXqqqWplGU0uHpy+hVhKq2dvH08T9M99ddKbRZNFL23bC83uutu2Yqc+qUTvvtOHxFj8Mt2
J0DnKLxtYYMZi3czN4H06Fb7sDbM6+vmZZKn+yv+PZXt0vCWmMEhxWCoItaBLGJXyPTMZwGi6Emx
FD2qOtakYnf5pDzSN1KSxgCAblJw/FlOzlROzqJAEFzf1SeUBV7fLgEPpreVq0dKXnUS4JBCewoQ
POW/fyiRVqCrf8rP3KBynJOuwUNh20AN355Og/4FH/jJjLn+XmtwPJVd57ekfSCjnvauEPiM146T
enNaRcrgAw26bus70Z6yKVA23fedYK2ZeyznnHDcmRBE6jZzW+cWx7BgdgK0rlQUPSRJwn/CecJ/
2bgQONF1GsXOFoaOno7AryucZUSufWu+LrPblQAs50PxW46nxz55V/W2D78jdygfQosaplKWzqco
J7R9bV+OMfk4bwlZfj3ynXQrAr0C+5pQxPErdp4JPN3oe8+IEo13EcVyvXWrwwH1U9sWtq2HjLs+
M4DlHkq+F18iBdtv6mN6Lb/BRLuu5ocm10fLV1W2iac+brdQNT609pCj+XYT1JCVbA3tSQyCiWY9
TXO1dNTrRuKWpwr3CcKk3MmkALUDDgE6R3+cOBHsw1R8+oGsy0rpZ1847x+mKwP8+xIB8eyCTa3f
8pIY97ZPE0OXd/5+r8rI4Xb/e1oHpv8L8xwquXtQ3swDOLy2Gbtqy72VnjfE2sv7ai0wAvdX7PG9
OeFyI0L9WM/C5C9t8X8ZLmEpOISfWgWID15elO70vV7gWzR1QWBuNwVFlERgVEyOVf8z1R7/rH9M
YglMYm4mL/hA5thj6qPEO4eK0bYdj7AlS97j0K0qUc/1vMWsgNCplYObtWPTjxsEOvksR3AJptd3
ugrUG9wpCq8+9JfsNEU4pIRBkCbKHxYNh+pyOUKyDvLn20LWZYMH0ZCYKt8D4D46nPmVUfAIrSrQ
wNxvfmKhy9XfuaDtsG9NGD8VgaAgTmpbcCzuZjl4fmRcTWqHDyGRmidXtW+20NmKnj+InYWoDSNC
VyU0gdoI3Is3p5dJYilY5aRJedFvP3jMCDCKI1gtYRw5m4mNEEn9yfa2iLUb6b5YQnzrt0nLfX5a
FAF0rKfZsmex0yGdsnqstlHtNySGCyF3N8N5/9vct6+SgV66xBYpo5bctBmhLcC62q6M99rmOz0f
tbosoyMzpYz4J3Gp7um85sIpVpzzg9qEsUY7LHgXhTOAL4CR/I9eUMH0mgjWvcPl+Ge6cAmX8kDx
SaqtlIVDj/rB/5CMZW09RsyKpJSbDSJ0Va+6I9V7zoAZtnVocIrQjGwrtSKHUm1uIBlQoC0kCd22
13UGto9aqar/RyrZEwpZE7KhYnFmtbaCzlSgK+f+5WhW3tue0TGaA+nmAJr81tbx5G1kOaypboaT
Y8olGf1c3Q4mtvFsOomKkczWsTzcxwlJf1030s37dlBq9bISJSc4fFw65XmBVMPwgGZQ0doTMwuu
YSfHxRliYIhl8wMbo59ozQytOr0KeNdXbI+ZQVLu7ExOTJAzt9iRhF8Qv9AZgOJHfqAZn2pVunOG
ioSYebmu+wvj9zildCV5Uhaw15Yx4Glc24tgxohktoue
`pragma protect end_protected
