module axi_wrapper(input a, output b);

endmodule