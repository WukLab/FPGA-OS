`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
HqZOgSldqG5tvTCRf1zs+dphl5cUc/CliJwNOzdNG01xo2LhuzjPfio7E4moyXOnUc3K822gOC2J
TYESLZa6Ew==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
OIrDoaKHbNNpNa4Y8RUB2UPr3sEL+El5NrG/WRqCn6FNNDoR4UzBLdZ0RkEtE/kd1e8qiRAXnNAS
ntmLbCfIDRGouwVdBI9quOd2c6niuf0l1ifPdNydgTlmdcvcH4FtGWwbj0s7XJFHWWMmUYrK7Oa7
ypoX0yI8X9ofX8I6gZE=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
o2BaFuqty9flAznx/M8gNeFxdG+6BtCsR2aqsQ/9DAHxxCg/poCm83GKW3D5l1CyH2rssJb6cxkk
Eu4wYCF3+WbM6vMZ9f+ue/D+d8YTYeFQkvn/1YGbQMdJFvnA7APNGpNaEdHyTA++bvpHcLeDHXmZ
UHcO2oKDRCktMQfkIpWYl5Uo5X9XXUuSCErwm4mO+pabJTx10qFJm+2t7GFI7XW8OT4n0wCvSYgY
saFw/TFIQDvcVztOh2fob5HQv+TFN1PaJ1d0pMPHd56zhCMoIK/tpXtc30Jq5rC3AYUlrAVI7rWh
xSej7spjHO8KQGW4glNrsKHlKmgtmQkDy5lgow==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
rmvJ2i95uwX6niiAKyEcn4w5a5jwqwFDSSCzkuRRPy5uADfO9kTtGpY9xAg4nH/sFUrTqV5N3YPq
0BdNKP6gSGLrEJkoXOootZZppHhpdq5iRFvBXvZxrgdCj2HjbkqgVI28QIB+y298YTDVRj5b68lk
3XM4djz0astyWqKuTfiHEQOzdAh4V2AWsKw90RWVDMwlohtbmSitOglZaKgt5Agn8PIuHUEmEy3C
ztCXVJSBJcg39swaCvjqJCetqH8sDtdnD9mIBT1HftWhwZE1e7lyikmHnfmfK8vuw4T33h5Gape7
vnnIgrdbZB2W2VQIABZt71DsxlxHEyiPboWV1w==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
FeRG0gFDBBAOsAnHq5GViJdFo6Qb1ZFT0UL3wMJxW4ftZOtVWkNDkaE5UmxGJJ0f9gF24avnN1ZL
d3QhmOmBoZ8JbNoIiI7J1MrlDHAbBN/ifpmT/b7LxeYXKOiCFQO/zFVofVLz21G6IsBvYupzS+Vd
LwgjRJmaalcUKVH4UosVym+/C2zusZ+Ak5Bm2dvaJGMhvy3dk0jKFBHj0FhAcguCB5muoY9GXeE6
qsi55D+yfO467kyfwF+C5abKRwtauELmOvL8F35igP+6aFoA6jkkJ9+n6dWupBWVNRdBXSI/OVFQ
kt3hdJO8GPFYe8pbdejonab7nXq1DSML+ln6nA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
FpxVfDEAB0B5LkPMMG5hGqu+hnzUCzZPbmR6wUNWvXUGjy5JMgXBybn5e1QSIgafyvSRQbfTya5d
NosrLSTzCxhpGOOURooEpIYzgAP9stuifgRqARx426tnZTAVojulCTnEH5xxRr1Mk1KK5PdfKzg+
1aFoC+E5ZIF7o3SKLpU=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
MM97qkj3XYJ6oP46XdiQ39lI7hpjEEvWojGHibvflKBlJjxpl+AxaCTIShChhd7ks8VAgtrP+MYB
Lqy5MryjVqFfWHfuIcqhfDUjuCZiwVSjiX12PNtS871/Zi4nLu+sVaMdP9FLpiY1QANhBpL+E7rs
r4DOOzhpulqpELeV3idwcc/l8RlHDNT5+OaiPA454UjnKcVMkKDe7cz5sloGMTTxAg72GQmayB8f
ech8lV6BwrAUh9fRB0PjZ7DYgcn0TrZUcZ7edpuaPxciUaJHC7BXmGgdu187qByspEX0sKPA7QnU
jhczJXNugjarg44QWZCsO/8QJiUKCQXMueCYkw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 15104)
`pragma protect data_block
0VBXmFbxdP5Mqca2eQZg18tnyKA3z5alyU2aLPXgyCkduCf2K9s9ZJt0MnEkCvZfN2ztrRTKTz/s
HEp9f+58awO2Xfqm8gMUipKz1q+0V5AFVMEgU3D2sGncalBsThChlRZNi1luAmBALjitrHBJ63oY
ES1JeQHkf1Ey1Gng5cYL9IrTcYiWIjurFx7Qz5vm4dtpcK8vQkDJH4CGB0d0kpEQ4egD2X+bgJjC
8gL8fiPccumOoPzmbtMD0g9SBjrp4rfS7pkJ/7l/mcXCa1v37iqbKpDMy3miKvQ0P1htXqZZJRLy
H+S0goA7zzXfDJX3LBbfOpns6Fg3N9nGWvPo1ASnqTNL9K9KqSP22YkanpViU/3prIDFbtMnbr9R
cU7DuAXN9BehmrZdB3rxNzruLLD7l/BDggP9yjlozAGipMJ2gB2ZVM+06lDiojpI4kecDGbEqDIv
ztdx7I6MCHNT9ZYyHmsoGWdgJEWQjfoOM0iJFbYCsK3hOfVSENjLnlP7ODPQbKJBdEjzz99POgKH
GHdg7gl1MLIdT1nXgukD5Mw+lQCzHF7ioNIjzWrfkpwmrF1+KzPZ71FIfCBpJb0YXaHhX2peGmHr
CFXI4JVWZQzocj+pixGZmcdLjznjSzWfnF67nxge9fHcL3wQgPcpkcYVBztXLmfGkrPrBytf4N0E
TeOH+cn1Ecs+j+jVmfhOS3fg+ZTjqrQuB4uY1lsykLfTRDVyfn7XzLTzK58lSdeIkl+EwHvBR13F
Y9t5rY8dcXIVobmzXvJLsmTxzU2Q7YMK5r2W7bGBheSx8s+0YvxxXLuWG2BRfjoD1Wo/jhWWzEE/
1cMDKJRaV/jsleJdRGX54Pu4MDO0zNysDL1uHoubp17TUgn5jZW7EH2/CdSRRDxO8rNWfhJsemoh
71IuUlIzekMXvBEuNS4ArTRczO+QXnKku/RsRi3I0xN9lyg1MaSGOZtiOmv/Z0fi99hwOneEwgsD
KGXMofIjRUKOvmeRJxOZil+Wg4TXbSdWIqi2gDN7DSoj7EFoNfBFAbgel+JEeLmEQJi+K1kwgsZw
ocg5cPaAR0zNDZoC13gfosK+kIGsFZbPloEOSayKy4ge2mkV0EwZj1ORoePdVetIPZHvbHeKf6zW
xcP2JGyE5jvGwbakVvEvqOjgS0tudPwC5bUlYXDaYKds64F/BnzrgNXhBXKemqKPo9fqxvN0r/Za
XOtFruJ4UAeiaKkha/nlEcTdgwbXAKxFTu7XIXYxpATIrINU1xf6vdBul7LWMKbRRMBhGW+ffzf8
/QavawhFjeoR/Ed0OH/a2K8bZoBi8SlhYL2eULuxOzJwHsLvSGwaw+zVaVEfOnaAktObEvM0xlAF
dattbx1XnRhWj4Rwk5kyzmQ+Ys2ICLOOYF1jJ/kmb4aPNhNZ0BgYINRP3y+YtPErHCMSBdEdA31g
GDQht4JWY+BJhlJNdhEC3sv+/rdXz7Dcb77Gr/sbLZy3XgeS8WRsYAXVcXzwvPF15XnDF5nDGQ/H
PblhJaJc6TiJki6ZO2vx30+7qg2SXlymTrL+LqcqVDev9JfxglNm+WqntNx6x5JtcgxqkaeWVk7y
FoMp49v4uxpRLrjOXh3ywCc3SUEyzI1RMnsLSTSMy+oQR9GpWZw539sfyuyyK0S8WIaH4HXJKuA5
75oh6hcDTtEiP2uCng0q3ZZr6yJqd++eCZijGN+YcVtKyDK29QgBX27D3+f8+xVV0cg2N8XKxv0c
jb85l0YtW2YZzmykFX2CmH8sWyw8Ox+NKFq5WYp7Yr+hf/isKal/6M1Mwp8OCNekUNqC0oBdYoFk
Win2zhw5zmj8Zy0+cVChnFKSJSVZQhedym3V3Bv9VoQ7cqphii6sHcxGmuKgPAlpXRhDpIkDKID9
Yinj3Ux2Xim2r3+2eyOXWnFK5AtSe1dqXlsRlnMhfzTUF14xHUODbrDDfSW4SyIfU8Cu3uEdI5U3
jS47eT+noFoTDM0gURyY+gZ7XtKPO/nqsm6CjZ79jwAI3jKpzCVPO/xri9KKTOdvSe/YFwlxzy54
HPPrCkgX0UigqpEi0xS8NgInN3p4i+fIW1LRGnEjhLX+GgzklV9VAsIaACBSncJz9+5QYf5NZci8
dHUlKtywnAi5iSWucY6ZTZ7BtmoMOh6tWHUCQLYVabzuG++wPR0KW+FE4hz5MV3PtnDYbM+3hcAL
2WB5csVz9dO1mgRxBufZJccMdWD7LWuYUVV1ilBnbfh+imXehKXH/x/Tbxsj+5U9l4BFavbbLBP1
ulSclXnh0OpwLgTZCSOHCJIvOmtXex8h838CPG8zZZAgA9hEzYywhbtA/APEDoj5FNKk5cTwiy8v
EjxtocMGUXDQkK8ZYbyhynwo4obpyjB2gqPMkidJvmVCtGadXaJoppGd6ZATmbI4YCVdH3P++1/c
KUIXrcRrDU5GY/alNbHlP/4I59VTqNwfQ++BnHzU/Sr1EEOYaT8TUZ7op1ghsPfEAmk1yodc7hXM
xIL66DjtZuTAM1YTa3UfMRwToUgZ7j8NI75TcrgwMWOGJ9lHL3/vqBcjF5IKa1HsAOUrGqXWXbCi
Sea2wm77GX6V7bE4xxIZLfVjesS68EUm6t2uiZwQXoTABElXbJWPRs6a2Nf7J9wJGoR9gV68mvpo
F60Suay2wQ9/Y5+MQxPfoKtc0+LG2ckQ1X+EazsHxAZbLjubJNq7dhPa4faLTDnaBvsgx5QCCNpb
YppDW1DGfdg2endiZkAuMWiSrRhE9yFfxV0cGAUob4rHV13XEZ2gI7JD7xIdwrS7RkSSsD09X2pR
ZEBekvW/15niowoI+rA1CGLrv1HYIPEhhxV5hut+ZjRpJ+9RSYpu7Mssi0XTkpLskc8Wi7klRoYB
BiCo0L+GuI6llNaSVKoWVzOB1Dcf1Co5F4ctkh5Yek3Tt37pImr3k7+UjN/tqRNHnSuMWrve0lDB
ZwUuH3wa73uLkX2wV0ZNMQF72VX3R+JOc7g7BVazsrgniT//P4/ziL28U30fYZzm71B5CUcF5IEc
JndbzssnUEzfNdrQliyRTrPDF3PsCr2ZiTvnvNgARpD59jtthAchDBs769y8xkFCc3dH5hdQjhJW
Uwzx/++nnc2pGbFo1vMXxCNF6rOkX/LCxrvx1ATgglwgwLIkh37r9ZXjV+5O8JZadXfxlI5Jth6J
9fvCPqjoNSKiplbq8kzy0V0WUe+JFWPHD2JOseOW/siIcr4+HgunWan8yWlwYdyLLcvSE650Sz90
eQaI20fzYvccgYdUTro1v0047xZX+Riwi0Ix6WC6Xml7v8S6s0gZ5vIZE8fUGjW8nhJKu1fFMErx
2LF8p2isVCZEMoAxPOqGDbM02QdmOZS8FIGJrN/zRv/UT4wR38i2jnJuWJO7NRFVR+fm56nYcsxI
mY8Quo4tfjdtBvvdazQDunRuziSXZ016JDwANz+lAwryj/WPVMR3wwtJvhJoL2uxxNy8Bj33MVLe
brRhuoeNlCq0DSmnhfcHvIIbwCfTcysfkHRxvrLzSIUNLVNS4jVaX1PlNaTeVw/Sq/Dp5pXeKKbV
NXdrB0+QtkwY2ahkM4vvM75loStm34ARLxNfVVIOwjWOEpiJLL7AbbHMNa+ukRgrtQbCKGVfm9P8
FmCkN+kzXMnjQ8M4BG46Iga6Y12FOa+2BaaEEcmDTD7OgDOIb67RQCrhRvCwEAdOg2eTXKhnTCql
WsGGDkc+CNDGzsxTEc66ZQavXGBSzra6R3+YTL2BNYeFijOd1rsucEsmVaVcrF0Q5LHnDjzce2ge
+G/zxurxUj/iym/sTYBpcqJ++rubM+oicq/SZbOXeoO+dNIQsZDyQXj5H9AFvepQ43TNCXZuaMfy
lKQEc5jiCijdMTb0VT9kIVknVgnOSD/KzLcRKim7oUV0T69YfyO9HxmL/Xd/Fbm34zLnUFMX3BRv
a4S6/ojIOvejuS4FZLoDQP/WBz9A2SbhR9LWe6Pn2WNsBznwEsKWAJvC3PtO/A0tmNdxpwZAcCwN
Mg9F//BEcsWcl8+bmsYM3MGlgKE54BjuYzZG7omIozAxlDELhPBERJ9PbOyzVTY/VWe4pg6fS4vT
REfDNWjZdwnggW2hbw8eYEDk2iyrhnr+nE4f36DwbjDuGYaDkOo4wt0b115emn9lNSWebcmiJY+l
ybTSlenbcoMMXChJDxl10Tvxo7rJwPJMQpKy/CwtANoMmQgt0pfomXIXGv7NO2YD2H2q/1uNJkFH
EQOCPadHYVFuJboK9eWE5Bg6s151XG+2Dt0Lfnl6GuxiwxFnn3UnEjQF5QeS7tZT2ANxVmHUrhgo
RvVlb6zKy68CXjmt+XhUmCjE7rRV1DqNTt1+m6H6b4XBx2ueSQ3hPRh1/cpDIzq8FUzS8QzKmcGk
tMxZHve6UyfsD3heDUzfafOQ32/q9HtPrHwsNrmsVzjPwk/enhyHrjhvNbewOwMNa0AkJIwxBbT1
jgdEq0/FC9FfwuQSMKBSEWBl4H4JYscRU2Q7hXwgfJe28q3gal9YbTk/Di+NIljbyLgxmU53ZMup
Xhuf/Ax23FUBI3ER+184wHDlR6z1dd6icGB+X77abY/S+5wCQRhWgDekJnt/PO3STOd8LUsE1MLw
SUOpqDwNnkEOye3ExCQE+IgYENnE6rsknIktRi05LQ/8IRvdLX1EP8CXry2XsNzyM4lvQyl6hrqv
F0lk3frQ86xjoKxq/H1VraikUhI5iP2D4Ze/JIiiA/DDSkIMQCqiRY/FLpigh0g2Xb375llBsnbg
+GOfI7mAFGTYKoMHRyRH+HRH18m5RtLk6LS2cTdVJuWj15Ywar18pOQinyC/sy1JrI7sK4P3/BIz
DTiIlxPIsliBfYThJuEqsVgTKfoBrmlbDbk7T6NfLCD4IbYgoLPghsyuI8ekk8ucXMcCUYzQRwcP
ERe53A1KkqO8haZpi8bOm6sCuNoptOR04ozaHx/F0k7TtwfoS1DTy0qtpTvmseKHJ9h2ndXfwKwV
jU3Q7h9hDIn0y1xSXiizPAf3wj6trJuesrQD8SLTv9b0zob/lnT8mxiS3rz3nptdCGmMjV9mj20E
Cte2bUNWq91Y7K5ygiNVVaVgFFQh5cZ/FVyxVdqjLasOYt4gVQCfaz/zps5leAR6Wde8WopqAXDf
QFP9w10Ebo6NvckTv0X/A4ES648f5wfAtBbii1u4iUSpBC4ELbuGG0hKkjsg0u0+Jzu7yiln10W1
tVNYfEPgJwZleiz3AIVlNEH4xtEM6AAyLu70koBl1717F9R6c2vjH90NPbNlhVQSap9zNCT8YRLr
6pn9OZibs8OkVyo3wNHLEHse/HDOa/KYNh5eSw64avWlysV+Gwd0JWgOzPfktBaVNL0aGqyaVrp7
yk1I09O5VnR6OUxZm67mwQ4BvHC6/fYY21kEpQbbLFJWQlruZGYaQF+S7p0fbW5SBQRK9KDwOg0/
iTOs09SdneXir5+1RQekKcvOxcEUWl9gTwzJhJ6HzH39uWW5u6XIpMsGL7NMQPu4ljWqqafm8v3j
3mahl9/uoM8V3I0JYmSMYKCjl9tVf/413RbgJT6e2GWAoxpDMVq1IA+C6MVM+nQXafQCe5BWz/JD
V3c5hOlWOdjSw/0l99vQaW5eVrnqdsNsZQYpZy2dkQTq6KOluy94KHwD8XO/yqeuR6CrMQeMUjJ7
vNVDY+5nTqn9Sjb4lzn4/UGq9JloN7mblmz8YtefrN572FViWJkjHWh4NQcX8/o9hm+gAeTnv6hP
N4/H/INTrhYhchUbGxpu5nP6r5u/gmdmPJQ4CgbiEko7cpAi5qx8kOxEQetLcrgpOXxX5dmu9EEk
rDlAlfC9bx1AU+DDKVoF9FzrdxzwYkPJAG3OAgEIdt264sF51uoDL/P/ApWJ8L4cy69CRoPYMF8j
4mt1QrV0uOx6l2a0oleVw7TwEdpSIOBHzqwEbxdtr5AVHVd6dwcATl73344nwmDlN5ROkBdfEHbu
Pji2lV5j4oj4tMPfG2n+groPpSJ4Z7bmNTtMnc+bhY66saFdfOdihBBrESDM0xG1Tjs1/p7h9a0h
cNRkzUv0Yj/BQ3HAN56lXXQmJnfyJAMnC3ZXtw/C8IIkWZk2G0asL0vzKJmK9LlrC8ZqkVikBQ9s
iT9YSamADvH9rZ4M4xoWnyKX5HtjzfxruVpuRjHOeCL2so6NPK/n3rFuyoMSEu0x+wlelIcJJ7lW
PuHjFo/HYHBGDh5lC2gwiUCIdP3U6gqR5tZRzrc+C/aZ6lyLniE3RGMnzzhEk5AIOf6s41FpGIKm
STc/D1IFWOzaba5bBhzhK/FAxOeLX1/o8ksd3R0d7PmDV0kFPgkiWn3gDDaeskgDhA+bwVf16HKb
rjX+mxrxvIPFVt5sxfhJbZUHsluW6gV1pwrFPBhcv7S5eWQrMruz7/fqrpklOh4gKL7cjqdxmgH9
WfreFBzB4OzxEiqAZs2qphR0O4p5vbAdXbJsRkXcG6nP3lm1N73RPL/zhblA7Dt/8CCt0F+M7ZM1
LYUYgExtmIZKLz96iQBzN3Top1C2/TyvVkO2QWpIo4TENdKa17c3FIzAFGs4UVEQIfj4obI4I+ET
d4aFOpoBBUPjBW+uPFcYjM9lV3z/iOsaXwKovnKZpHE5zYlub21G+UcmEC8KG6ghc0MW65/vATPS
kGMryd58wrPE5MY3RxteSs3YSKXM33xCD0w8EQPhCyUXtMnWlVFtNmMSVLGW2ZWJQP2QJWzkuYW3
6nZB7yBaIHiA98hYrHQy+KE0b8CqHWCOYT6ZbrRPpRywuQoN8ad3Cp2ZLRplQd0pHQ0dBiN0imYP
TtBIzyZdoWoMCil3hN61zIISF3VXnicKT9+1upkE2JjnEcuCNzHd5Uwnht+i037jUoVsi+wdatW8
vFiVXOZ4DDrLSNbJ7rjT2V6uak8w7p6hrqhoUVdvvLhZvFQbEv/j5Y6E+Zu6blu9WRJYvjwSjvjq
Jm5ukFjVqAv7tIdrO47shnyGjs5dKo/4kb5ElHAdddZC1c1WKuju6rw5WDDS/0p9l74HxCgis+sf
YTL5XAZp8Ywjl4xrXlvEWna+9RA1kAD2V71vin9UQAE7yUUf8aMbMOpvxDYpSbs6C7Hi5koPiZ1t
5jinDvcPPF+st/cN2ruyQkKCNVMREBqESk/wWLpx5TzOxjtv0jB7m31N0ycTj4E+uya7dhI364Sm
BeLDUDe2M/2MJDsCZp034AvmQjPSdww6m7wpOqLf5ylRwYw+MiIODq56p/wzxFwC7VCeg7hxz+GL
h6+wSceLjhCQISvmXqNONp9gR6WxkS+NCEpG6bxRL6rY/PAFicYuUXAXCNQzFMjLTweW6BdkK8qF
cc7/q7y0JPcEHHXLlhV4uvBWYlyaPdMLm3f2Q6BWXbfiSaultQRNrYI49iM8Z6WP69G74Pla4G55
yxasWlB+bOlmGMcOd7XV0Q/0hFSKaXok0RB4FHQqReY49/uAV4bQ+sejHz6i8ppXR/gYyZaB8UZM
7lgnEBJO5zDSbuzsgDxfcE0bY2TKv66iLrTjcyOET+oyPrBHLN44M609BXKUkp9d4yjETAkgCVba
/UYN+tUA3/UcwdK9y4HCDpjtiUUw1Rx3kJYMyIrxnlldqkf1+CQmw5PY26cG0xYs5HD1j8mJfrBh
WrXRYL5Dhvv3s8HzVYJDbgOHPCAdPsi50AWFGhDFwdWUXzEL3h7sWAwqEPuP6kPZBc0O3ACgkxls
vl5ggSlR2R6s+i0yKI5I21DhgvYGsMIsXerRUYrABC8XRXC56EVYDkgK0q5mQkrkT7K589KrXh1+
yWoI7oCTKwX65qCuHsBAxmr+UlMLXrAZ/6YDE2Z3x7lcEpa/y0VxhgEetBs7kf2bT93f1dTXRRy7
cH04Y79pwMxSc9bk+147VGM1URYMqKdIVhUFtw4TohdQyQYj4/xoSQlCmdUO3Sc6+AqGW8PMiKHF
jcIwj5dlumnhvEQGSX9bY7VY5qu3Qnsg+pmuUl9qzWGLM47X0Z2epTYbTZ6fY7QYf7iew5OPg2Zf
cu1n6DItdgpGWRFp3VCvC8LMJC/6AOxYKpPgYX5Ji/yHcwyLGXTAxdxz0yltm1yWXvNxdYyTDpxJ
KYlgRgBogZHhcSA+OrpBE4OgKWhRGpuGR2o2NJwkGzIXPba/vsK9SmaeF/1+E6h+AqKFxrVIGRb2
OgY56FgZHTPfyPB2czuZXFhS7UKQEkbkl8y5C483BseWuy2sTRoAqL9sNDOIlDQKwkcxsyQeJekD
+dGAalJaec5LuHj4SbySg9cGFleRS3I21H62/tbt6yappKI+wjRnp80xEyIg2nx37GcG5SA30Y39
gKWM6f1c1HJDh9BJZrn2aQlctlggk8ugN1kJadhdgMQkSv/WT8BAZJRsXaWUTx4si22UmqMESMh0
dHMvSAfkVUtYvpuW5ZWsbCmWMFZaLGpK6jq+qO3gCOgKhNQJLFEEuiQYvqY+rbaoi1GppycrCNzY
pJDsa73JZ6AvmaeLju9IKR0TKdQlDgGTZm6GhVVFQxLB8qAjSdnjaIceEAMiUZjqWBAnV6C8xJhP
P7PduzBlHegw8TvPul74vP89BztIuP/Bm24FJO5k+RKKZY7IFpAJ32zAc+PYBPmpQY5Du94tVXhH
V+l7YJMdL3syuCgKtxur3aQxr2RzfWBgzmPvfdIxvx9zknWzV1tsF3Zas8s08q7pSLNt7+UlDW7w
Ue8n4PWfeapHVwMMfh+ak8C9nDYwP9KfscGDUmG58pt4Y0XHRiBibYId6ns+4vva5Ua8qB4Sy1jY
u31k7BiDGakJ3Y/DBJE1eO+Z58Nea4+jJ4Ke1Z38DRPVJbCWzhvtPznmmvOSaaceJkEV6A8G1Ivo
P4PIs33JdGFkw0wjeOcK+dVZfz1XiiAzxn7qUvQvDWqjKJqeF7OgzR5FyIRGXifzl3k+2ygwtABl
Bmtsj2s2K67MqrI6n8XgriVbR28ARtv6zJ6riFrDqoRIVkwXCepnmghwYC0xk1NQHKJxOjQHAEZA
RpQwrPzthG8FqhSN+YgmT28SY4ZOnnvQILVkUwsCU1P+S23aam9kCubfpo5tDvuvIDVCk7Kd7ECs
jJIWVsPhu9IOrfsc444yWFugVbgdMSGK6f9WBr9FjCGgS/N36mcREHX32vlZ+5QvgvkZ1xrqVx2D
n63U7EAoZUHnQDkh1o/0Xza0JXM4cmcdPDdymsSI51QK8NVUY41Nzgh0E/WxKk0wkCsBl6RLowYV
SSK6MMW7nkkefzBSgEBgz7CuI3EdWA20vkll3Wujuib9nqrl4fGd1ArxaP4KlKqHMuRX6sertDTm
FkEo8DtBzxd3eAHR2UX6fvXqRcKRBd8DknLHELhlTcbwqCpmtBjW9WHAbDadkJWCl5o9Wd1goR0p
ar7a7Vaj2kMJ8AVMEQQ/mbGvI6ioIik+MjEY0rjm+0fIWTNbII4v356R7aT5FgPOoEeuVRWIvLZy
X10HphrlYa9i4Z/Hbvp2x1ygzy7FwuOQi0rdAbhOg5+z1NG+0TfxihfgDETL5pISL/W61+hrar8b
2s4njvJvHuq5zKp4R9IPn6g6T3NmhgvmMNUWkA3THjr5O5oI+k577f/kavaxxV/BbPmAlK6aokFy
QX5zE4wGntsyJXVf/4tNKYpt8bnBv2KCsFkpVjj1NUFcX1bsoOsCmjtibBqMSDzEniMrH7cEMSK5
T8Wk28vmncY0o8vvuB6Fz4TfeRsvos87Wz3JHoC3B3ATPVRzEWEhE3lcxyVl3Z+vdUqIzoIp42Qg
8iLFoMZVl7zLdFTGm5LTn1yeXJ03/lBfBjUyI0/XsmOahchPytyJJJjy4v7iCVkl1VBrIYUaRW0s
1+SlhZJXTTJuS8IOoWDAmKMj+k6LXre9o9/kOL+6Kw5K1wHCnGifFXXW3h7NR9tLpQgQ+pdaps5O
z+eN3Rf+eSb4e9ZGB8Dfrehk8sVqywSsdy9qmZjs9Geeh0GySfvfoJ/pMG9ibugot8ma+34E1r6Z
4DxH6RKM9MU39BUTmuPsyMXAdo13P8PIw/7Q+JzSFVK3M83btC5xpismCDH7BRtExQGNrhaBf3hy
kjMTciQ1wODaHDpfRE0P2DNJZOhfQeJTNhBIMAkSjV2/iRIkpIMOkYmh2CSBbJ7xrYC1LAtmC2W0
TmEh5ljuPPqIzgL7GDBUmFO02/mCq0h2/b/bOeKw0jnLr+nAiznXD2hQvhbe8aeszGxXpU4RZmvo
4L8QFpBM9jEs+819jkH12VUNY99PWQfIAATQIPFQxByLQRPmrkVPbDI7vfAzsxYcdDHVZTbG1kRZ
fhobUKxHWcdmvoKHbgMzczzOUXgb+b2+CV8mgt1uz6dIvur8Noi2wIgDiSxgLnWm0d0PDiSZsI9N
RkCaeh6uwF65ydrvgzmTLgNtCfi3Y6+WKz8WxTq1wt+UAYs1nMnFVZo095kue2DHMMQtUvBaiwNn
lndvMoNiFvRbuqqQVpri3pUotJnVHUAuClTCpstx7SuphGOY5MbxZ2+JvAm9a3BdSrIpNoOW7eBY
OFyStl6dFzP88pL7OjEdVBoh+r8sRUVok1koYqcG04gzkkd8Qg4xOQtxc2y5hA0+5wNziqDEpo+z
yTOre0UxhSjIvZ2LYpcspkeiH2kpsawYdAxjdFh4jULDkqmj46nut2Utzz7zgmeEP6u4dV7M61n8
p59M4jQQ7GqzsqK+Ul4XY0sLqkp+W9AAWKd6szmlxdky6M/KRV891y+JZhPosL4J/u6NPqUDqx3e
Oqre/do+E3Xjqimj/eE4lUAnYtqCs/Y1BH7cFKVa3OmFuIt0HhRVnpBOOgShkDrCxT37UXhHqx8P
rGzsgpovrLGoeSbw1zABzjmj4OOl8ecUCy6vJEF3z+/wPrlKMtXsrZEfJpAWtiuz+qFEEm1MKxDs
Bf7hIOSKwWz2mlLrIFh+k8ex/RijBvTMg9f+OahoPb+8mMYH0608Ikttd5Cuh5ohsEc6L2lxIOWn
1hpz8e8Oulh9DECTvQ3/UlvUiFgmU6qHT0LeISLbx4O0ACjFInMKFKswloCNO4901j6n2mQfvdwD
tF2eBMIfYidvWjKrCSiYSW3eaMuGWQh0V7wjZiKpFLOkw0jddf3rMZC7B3fYVwRVW/Mt2nC59FmN
jFaaQjUkXbwYpZd20O59Z5JXZqGAgRDHHICC7EYKfP+4Jv662VE+4LfqanIpwUrwGj8thDVeF4kx
flMe58qBpDeEyy9gBW/XK2xpxN5gaBSQ91Qzg5NxOBrVVO523Yps+u9Cutg7tZDHNCia9kLXfmw5
o8sn8LtuqkZgES4aLGij95Dm6e1EkklYipmkdaVEHh+PUTlOT4AdqgxM+RZJZV5tuedmYsKYSNsG
hdxYNMHTt46p7ftwqo97yIhvHC2WGAzVvn/RzXPWdZ2wxwmYfUvCIQtvpV/6fogCZqwCVSO0HTDF
bqx9R+PFqlUFiqCesHkGSWOmAtkqH1qPjaqEcLF2HbJHXpQrgDxbzEGceAm1m0vZLmnHSjk7OHVr
is9OikJp39ydcqJE6t5E8UNthcfd0DQOunxTUlnd3KXCVuodW7zddirPUIG6RlYtUnak6W/vQUdE
8EsjYA9R/U6pcpHJTIk+MApM4CwAcdiimph4KpM1MWZ3QwipWU5Y0mCQ2IRzTJL3/QA0/DqaTldC
xgKbhFi/jW7fb7SGFxSLjOrNxvvgQc8tQngnpXzqYWjmXgntgAtwFv4RwMm6RQ8D2ImLz6cOv051
wWzc2375fbcMKNaJ+PV4cm6SYGqaDaWuYw7lgTQDh4l3Y5RWJvjJeO1LhX/fqFu8w8Vs9Ev/EKV/
wI2y0oPC8eiiz8FQjU20rTo+z1sw6h8MM9StF5jcbDEsCUQwz3dVyj+zqzU3puyBRdT4K/88wjxa
sMzkEwXARorH60/5kGR/9L7CjlE+ibw0d9T5uBnH/U30PZp2HDZ2IcrEltEIRgeBdhNbFCTcrIf4
LRFDCxXZeNDr5SMnMrZTbB4I6uOv7oO5Mvwk/VwEjSFimJ6W3qyE+CJTwcYN5dGaWXdB4LDu1nYj
Ju+oqewkND5vwuta92XRUbmbP0N/xq0AjddOJSVlgsxsLZPrL2n0+l4Cl+CQioVgwrIpk/RxxJH3
yGTwz55a4vpt3slFRhwdTKC0NeqdNYuw1TRnW78wEkvNwAOlrse++gMNpY9LPv+J9db7MT3sLBAq
7Im4tFS+8Ll5GBXoTA7tcSbEKe5CM+1+Ha/Ci+/aLEmzzgwMsbwTnMsIEQHu0qbsMPrjranXJPFQ
IggylNkt9jOvA8SFP+YoPX5z8W1R7DKHaT8xLiE2AsTk0t3Y//9ljxKLyXqd31XGBi6z/Zqtc7fN
evekI3Mpk5Cfpd9oK7ga7pSni9GGnr3L9DacsIgiZqiLariqRX1hPnhY1peRAWDns9mddi+qm9xE
XzozNS2NhsRprHK6U9ulOCejPaRzv478/Hx9ob/GNWWMqsXmGs3jJREbLtxqrvV8ZrRs4NIOmOQy
bgiJSUCWklCEWs6ZzxCEwkgo8LbA/QyhQfmxMx9a4ji3KKjFV9GtTTIoMcZYmjU4FDUw0496iVK6
DmuD/VUiZwKKLOCO3r/mOpj/wbcoHDV8uc+453rvxmHyPg85fp/umIi2Uc2j5f/sGSx4lumZv4hR
9bNp8QaUG47gGSI5FO6AACg3fc0VQGsNeVg8BKC3dM4qK9AEbQOtquCExhD6OoKidE3zrNHcFB3f
kY8rnpU3yvRXfq4SLIbzcp5IWG2pv9zjsUI7LbIYu7azwOeLwX42hn4e6tpRsiOZ5BYlxm0pl+k8
qHnQWzyrJNECJevnHbygLu+/uCH1jI6xwPpnAMfTNnrswilDppwKlnE1/h4jxi+9Cgbjy/aOKYeu
d/iki3nQ/YMBHrbxNd1B0cDIYGlDpYDY6t19oohKjIqo4s9jDBXEFsZf+n1OLRznwIJnS4vlqzt4
cSsVeLKWluBitTr59cOPXZddyNB0aP7d0vebGEM49rdBhD9GKzcgrzwd7w/ljm/ITar5yzEoiMHM
YmeQA2T3jJA+Pbhy+73bowqdgpH7UUtkBRQZgom+ERgZKOPNNdOQk6eJyGskTHkanEi2HbdoWvy1
iyIo7TSQvwB4KqnaHJIBvTVbWmF62U2/nKq7rPTwwKP4DkHyWvf0ApwW4Qrng4OvQ4YweUM3CCZC
k16+NImcfG60YPJU6NCOIqM4AiuS2VBab3C+8PkbU6ycBaQh6HJyGCr57zktkq1OEZE6eKzXuKpI
2zpWCDqY1KKH5s0vmaZIAKvizUOFWpM18MsruNIUFSjhctfIiYnEq9CE2+4YBb5pnEsudyN3NSHg
hNqi81IEm3OQRWtiSLakVUjTy3bkXOXRSs5+7lqCVsGT2PPlNkW7EyYJb0OereAT4+8hyBrxcQpJ
AHHc/yORgc+j3o2iG+gD8KI3q5jASWi+nlr+hnX79DNZAX8W+Fjl96RpaFwenwQIDw9HRA3CVCU0
izpoh8Tnep89HRGTaL4zdlq46eq9+tOd8eOOTw7Tq9tLeWrr9D2KSUwkXgZ+iPY4kUoKKYNgqRdD
visCZ3JncHBe9eSxY5Qox17HhHo84oc/yF2sQLxcgZmj1kGfEt7eBtpm1l2zOTOTF3TvCe657pvv
OG5wcCgYGGsyF6TaxDDbn0dz8yk8ufbltEWYdJjXgr4I69FLpnyW6q1fmyVnVIx36H479w0rZn1b
YMA8mL5670QbQaHTGZHR79BVo7RCzdbtyb8JmwQVRRb44wGLBWx5JM0kMKKjKRpTj+SZ4H05mz+v
P/gBQSXePzyWpQj3YPMwrCrVR/hQT63K4S3jN4FiFI8R+y2gjA4yzKZuaxYzD/ywkVv8uCE1J7QF
2Deb1lg3BFI3SEy6Kmp6Hj8NNOfPLk/h7VXXrPGU2UhW55u5wwbG7edDQnvHKTPFjE6z50GALgai
6tX0WAj5XMG7I5LWBjnfwQ+L9llHDS8fDDLpAT7pfMvtImAPV58IaD4piFpPXeWL48/G5bd5xcdb
in9DyC9q95JvDtBETpHqFVBkNQI+Sedf6663Yostmbh8IVNTxOrUtTfUK2sWBPYfCTyNlEnq5+kH
S9cxrSYxNbnC+HJPbQaJC3v4+Wd1VMg8sFsSUjb+ykhsO8IL6qHLTaQD5Q+q6qa/xYzQgoGFInK0
49MQ+c29bwYkJK2lD3TtjMd2r8gIXBlpeM7lDMYP5zZJKobI9CILyTtNztvnzu3icY8Cg8YpVbsX
5A3/o42CO5A5I//srA4ME6/sabIYrY696BJ8vO22l96jbU4c+W2rN9N3ucp4oWxPLnGZMJvTmrHJ
hxf1LuSWvmpdkOEMXlE3DdwN7LzudyEBrXhn7f9sHPOVub2Qz3exz+x6+INVzIeEKQVQ/e9Dgh/n
8OIb9IMkWMaJ6DWfRUW7klPqoEtZMS1uJwgOzKLrbe07XZltWR5ne7LTAg/gz2j8lNIx1z0SzB7l
hjUrpSp1B6UKzORnFDVNT3nAYfYubLy+o1bxnVHbEL15LzbJ2qQERTm/pAwcUJgQB2PVoJhkYrZc
SsiuzMa/EyvfMZNmuNX6XbTsBaijiXz1aDNrfnH84cN/evTCmnPsqeQkcFUOD8ZGC4IJJF3RZBuE
f+2IARydKr2CYtBOJkq/fy2OKjm+IxPZXYMncaGEkQlIGifzgr6aUZhowAl9oWC8ImrmvK6PYFZY
VDnqC0RaJbHN3Qc2yuXYuIh2ESJpW1/kSC2Xjf5ggaCHtxg3qjOnk2p9HWKU85oYYMKfTzs7KpRB
mCdaVPOWHYbt0ZP7uIpAgylS7+1Pk096Q4Wl2PwBaFFC+42yrULC3SfX6aPrYQxc9AckpSemKSnQ
R1cHmy4yHZQErjYrmfEX/fXjRG7xAKkN3RUDzDr2djwlVstn5ybjEKqHOhQ3JzTAJ5ekcgS9iudX
BJwb226ALVB+kXb9N3/AGzN5N6CcTDGQ5Zo9BW/pkD3KH+nFRnMGrrxI0LWDdwZYu+bORjwjgFh/
9dVdiSpKFCQQ2MxuH52+Kgh9gXhDJiqXuDZdt3zpt+5oreH2cL8fOu///yMrAIW+Wf5gbZDDL5ZW
n3KN1BnqkJLV/KKorxIUXPas1u+Ym5vhHDCs4tYoRVo7lxMjcLPXMy24tF6fkAiNH8CyzDhVCSQm
Cod1riNw8Ab1eK6gpn8uxGHTdhXiRjI8nwJDqv+Sy1WgQKSGcJFo+3BlBKr2QANwTMyVtHBmE0Io
Py5qCnzxtijvkq6DJ5Nthl4PSzmJXCl4lloLZWcivVE5mQBSuZZDVRRweSzoHq/Xpiy8XMaPJiM/
qhsuhqNkPgw1y7J8Phtg5Gz76m6hxJfCjsf9nzV5vCy/UM1mLFdwZ6DG4/36yADCngfEvrSjTvPx
GKqrLbyc/N/V6GA/Qjf2kCBrtn8KeQeeGM33ygE0KgVVy0Gs4g7tAg4fJJGnJRWAeGhRmgLgCBXB
J9kOr0k2JD51jhdl6HLxCLWnpW1mNaMttFO/8lfxYE8+r+Xp4ZDMu0WcAagEGbKe5EG1kKFUsaam
riUam9oewgEiHoED9N0sWAz9i1wLudiaQu9PlLIISG2DDpvn8iZLtcgqv1H1x8YH93E4mBD0gLMR
TKOEvqMFab7Snb5eWeu1QeNF/cdhds8pUJrDUtZJe2izm6pSrr5nXEE5opePcNSKiN4yvIBafN+B
92qfYhAfFFv9jzpF357I5NNVUf8TXgqauOAJ5Ub919YecOsIormazXQFvZLLHsnverMrJ6ZOaXo4
GFrX4Z1Tl+kF0eg3uYM+3p6ilqQe1mkA3og3etbFajSiKgK68SdGISBKVM1WPnPeXDMAylu5JuxJ
0mxcPlraJjbjXX6b0I6bKUbCpkMeOch3NtUkc3Bc41H8Dy0oSc1mvU0t072iDJMHeSCRXfZTmaOR
Q8iVVZcmNx6KjxKR/+RDcQfmKP5OfGxdhRDFEOureYg7O0Hm3Q5PHTBk6v3h7vKqJsfGGw6sIZ0U
R7olaxUDuksvZ9CHGjd5WhPVqhr/AHlvjetFtLAIK3oNqw4K8kIe5Mkh2uFNtPi7oLBlNfI+kH5T
iSx/BZvIIgBailRhGgHiz0fk9cBHQe8OhUNwJZ30IE+dnlKrMW1KR5xi480w6uFnHe+igG4e1Vny
y77b11lgNMZP5IJ9eqQX+enyNek6ax667QcBqw9JSTG3vUI3O4/X5DeOan6+jIAL66X0n+tR8Dmx
JdoPLa9ke7oavlR7ko+OkD9QDGt3HN2Vke56+uTuKnJjHH1ZtFYUs4RpWgWb6WhB6COMVSEBTEqR
PUBzBGvOWNN+jmH7m7kLyPZX7xaMum5U44IhCrrNNwmEr6CgsvWwxpC92pSRW1l13SuvIcdpiMUf
3lRu6eWWcxEVo+njzyi+d2qhI5H3zyy9ydh+GsHvIZ1QUarydaf68FCHOUM+mMEIifiqU3F8v1Y7
9fxTvhs7LOigsb+EKFkPnxe+bXhFW7v1UNuqDlB4BVQhycezpgSpFkCvHYGEArZfT18co7Ui+Rq8
HCzSPdTCiz8hSzMODncjyYJ8drnP1/fZdXXgen72/ZPE2uHBPSaaeSclNiU05JBN4Bfl9sjpAr2k
GLCC5AiaM3U3Ahv94HO6F7pVqK1z4D0yZBMIUvt/n0lrn3PZh7lQsCYqRBOId8PwXkrMjCcBgFWX
gGnFYEQbOZTfmEmTOpYCgRgrXs26+zPRKaeGvOnhz8bG119v1hl1DRyVqlfCJ14tQuNXJUZSbHIV
W8+ceHsq/Q2NpZaJrpxaeUOVrsaoflV1Cl81Je2POJWyBvD4g52l+5UDw+TwJm+25kQZSJ42h3+O
pLtMbJiqDaRuUyKmCu8mpOx5QN/qeoelFX6sPQqQNZ+wT0MkUnaqwkEYyTA/lTOejjSvnvzA4Ay6
47j0LI7FhNGvMDX3zDrwIt6a7Rj7pCwHXIXy5oheP4czaBbinoIquFPjBrcOaMVDiSBYPLACyXu1
jjgkeOwrmecDGr9XM4j9YgNNS8lTVt9Pn+z68NH4X+1+miHlfltMHJKNj/qQ1jHfw8Wh8ab+bDjk
+rlVvs2VlxhLWKQlaIkiQoMU0K7Y8TwVWIXPyJ4EWL0jpvOP+bovrXTtBLrOWh/o/SXg9F44Vhwy
pGbOC/6GQNc3HELpQIbF5lQGD8T7VmcEKs3eRq6IhyBRSNNrtwYHkqzoGV/mgHRJRj+l6B/23RuF
4QHjXFCyvGKx5RLpH22g91+exEQhHxdXGzK4plfzGXzv8UaEUW+Db+ZQ0dp6ObWLE1veMKXKEASL
BS+8hx3MWK0Os22IO4+4hTrUCATRTXjQFLXq83xTmU1JrGMm6mkC+OYXnlD2GbVlN3Xq3yV/3KFw
GTnnDZRsEnMmu2bycQeX2Jmjkug7CTKrEmXt2MwC0tQyjBu4rkJb1myAQOidLdJFypbRIOjN3RHD
Tvp1vhh1kPeyZpz9vOPaKpTFAvWBsUydEOk6vkuUe6YHGQuSjJP94HRNfo3ithi9f8jYsTe82a71
+C9t0SfSM03g1+kGgRNQxXD+9XN7DYqV5Yl0sgPvNuzP7wm9hWI/iG4Y8p+var3lsdble+UA8Ymv
cWfFyQx49F8adczlUlEIlj+d37K3JFKK4I8F4Sytlkrk8Lg+09MNzJcqWPDwXxz/QH3XveHxXg5T
+cDKa/PAcDPKL5bT93T5EMUXlxBlAKlhAs9hiqJU/yro4ovRISaKGVOEESLc7V///yRklJE0glMR
JkEmd3jE0cyuUDfOPmqx+mnrVV2aw1iXuGNjg2878QeqVM0J2rSQdqkjHrTrLN3GTsHpcOZIXyrT
+MJwOer31gQxhz46+CFZPU9AngehWKjo8jqXv+dmkB68Yz3CJ9FePn6sxaw9N+IgzUv9Rt+DAwdE
YIKH7+lM0kTkyxKNyjKdZ7QXkWB+56KjJvABVkykDEX4HIHj9oVtWpIax2rrY5Y5f838yvktgOge
RuR4k+C2t/WqC897ThZU1tyhEtjSNso1ScRkA0mP2alffy+KQQ93AI6Q57kkci2nqN16z7MGS+96
I3UYznu8yMb1p5b/t7JkdacINdn0n9XVpVN7u4Y0rmAZwQEW6r1Va3T+0WO9kvOr5mTQOAVatwRn
X4UyYlnLZT6956SiLavqq1Ode3mu52c0M0jRgxyxYXbE2oJGjS5LQH4NsBrsHtNsGpBq3XeefMbK
klwvLgV1iH/voqFeyK8OF/YErVlHb0H8kZVhUNTDkTDmAkQ7QhFgSv7oJtzfpoT8evuiGl+LX2Dy
2CyV2phyXbcGgvQ5jp1j/mSSOW1JRksrAay4VSnIVSGvnKgH+eu6Xc6zG3xj7Am/MyTJingKSqHx
T+gnOA5fIPqDka2G7YXMIb9fb4slgx8l9EtSuZISpXRtnOzf6y0Ttyj0o1rZvmoWMzuCHFGQnKIW
igZjr83oT2tlnXgo377w/X+uIKX9uMn7Pn4/B2GEEIl+wZQzPPh/8f484SUOYOxe9035qjBphJkb
QhSCDvP9UipOUmgNIxR+HcmrSK0ifHZK0vP5H9CFeDLftLinPZT0a98+R4ssVJ9rESdEvb5Q8bkJ
RcdnCBgnqKoZHQyzGGNEw0dGHue59h+JzmM0ko+jx8Ez91dsxrkhcASLzCbDRPAj/KLngfR+0K0w
+u0tVfQqusPa382dvle6dCDqTv3PoZfEaU54xLoX87QqE/GbQq2NCutpwXWcmHI9R9j2l3aCuopw
OA3KXDKm01OWxSsUPrxGhpEuuclGIla665hgZWVmw6rEz5Oz52ZFYqLHyi3yqF+nxEQ4jgCqtWAF
3vrzUwX/QGOCoBlnscb2jvKRXJl8MyQyKbDP5Fxy/tSetKDC1eOZ3AYvahIaMN0W8dFDsS1pp5/I
16ytjUc9je5vFp7lwdWxTpU9Rh8Fauhx8MGBc9Agq5tdlpK39iQCg2RM08JF5XkGMJxLn2v/BMWc
5MOF/VkrzMzqXo25yJAcsehohJW6zxL54n3Xzt5PK5gR9F6IWCNHJDWxhuk7wqNXh+zSXIto6K4V
20s/pfHP9uIlv8kHPUAft5rbzgp6NOl+e4zlK5L1rMMYORQzZuXJC6oq8AsWdgUJv+iHJweA3xL2
xADfDnLUOdQpPagPBy7xSIgiBzkCttFIu0J0OaMQLNK6CGGAm7N9zJIPgG5rqDzKVhxacWPp+wR3
F8+V1eipKpVR8hJzcagE1IaZVH5DNxVMexH2JR9WUCWGLL2knJezWREpPmU09Iep1+J/JhBzapbC
jG63/5UmeK+9uktUqMMMwgj5o6teY6aeFsHBBwSwibu68lsjsvYBNXW+Vpjdrba8NqAYvuGE38eN
UQYpk60vu7wnm4fVCKFSrAUjs+ZfM3Xp8rKIOChf8i6m1QIFiHEYqApj0W/X+H5ZUTz8gMpC6nWu
cbEx8pGuhbvU8VZHJ7YmWUUSW5KzTflppoebtD/2CaNWseDRK6cVK6gbfBvmWGG9xQJxhcp/JbtZ
DpwtnvpD6qoAgPkMz5UXv+XtDH3mLYdBYby6ktqQAXFRgOsm7XMbLH1XDrfVqYrR2R4UJVNf81uU
jJUWKhwPPwJ3xXVJFjLMRZoZa7yeQIgUaoNUz+8PalLey2lb4BfmTO8kjWHSTanq63dNtCxhkSl1
feUErYPxf/iI1egV+6U9Q/PyLK9lLw6aGh6iRjFMmVqHsQnWX6nN8hjgyHAdLyM/qjfuKzclMNRH
5OZBdBtwaWROpFV1w9Te8TnzxDA5/qDOHuwS56QFGOunpCZ5uJB5JPc2OaCpSRI3d/rfnH632YUc
U/rWl3BSr43HWikDa6ULsJNH5a1nC5uTpmDlGvUtMMRr4yYiGf9lwX8cphNnuTJhLd9g2tKR+/Qt
2i2vlKsza/aWptf9k6VtvvI5a43+5yG46peyVq2Z43BNgG7sU/zKJi9Ee1xGHjEKNaJxM574ZLZW
Fcwh+OJ/ktTsq7aUKgyELyWGTPh2NQc2jGK3EUwHPrqAnEwEhKSAIdpvJWsMQX3X6FcDVYBm6vCH
NMA2So4SOgTGsESxi4T7On0NVKfEU/5jzDEJF+M1kzcFIgGpSByqvyxSlGxhwzK/qE9jN0Fy0XA=
`pragma protect end_protected
