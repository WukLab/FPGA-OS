`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
qD05XqEbILxNx1j2uIatkH/z4lBMJYJPU3OkDTHP7fz0wAmPHzR3Z3+USZlABhJoZ4BTMNcxeNPB
A/nUMCo+Cw==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
NlnI9DvqPNHZHFaUCDlTvLlvMs/V6VqLMjYnixZVN72ynK4uR2OfDXbrJK0EHTxVU9nOtl3wRAGO
gtbOSPgC1PcIa2x4XGAUaVC4tGx1DBpodcXz3r4/mdd+HyDoJSAe9JnAXPLMPAneLqXfKekg7Eix
GWsDA3y4ss1cUkzjxSM=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
D90vB50uHGcywYnCyqeEJuDy0uYBWdZWQXx+QsKCYcnDOiyUi2Gh6dA9GY39EkKtMJloUqK57aPo
t7+JB+bjuR6ihQOUPEgVY/Wf9w63+J/Ij4ZB5iXpadMTbU+bE9j+xG3rZCvi36agnId+XrigTKAJ
aOjHNZh/BzJX27N+Zfj2OLkLpUQjhjZWTofXth4qa+q2m8yDFHITS+KM554dmKZlY8Zwz+foQA/t
Sd6VnHLrUChxMT7nK9QoSIYM1+i3Lv9nwykdyeBf/0T+T+ESDfLw+9+vagZsIe1AqS4RcGy75Cmy
Hq9aDJM5zGZ59KlgnY5jzQ9/K2MfiQBPufCBcQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
TX6g1Fc+0882cOzX3jthos5j2q5ZMbjsgs+KF+BMWBQH+QNYKtGT2oDBSMF3fsOPTql3jYVaO2Uc
yntwVuoX15AXuRq27aMAxkmleJzmRxC0ghbJ1GFb1BTl6Xe7vK+U47p6TmZrDUJ6JYG3KwGwW3wk
EYIPi9kyM3rqpSRRTyrlvBh/isgX3A7iUe/BpC0Jj+y+XyJYckiUoyPttJpPcEb4egG3mAvoWjnN
70gpIqXoctHuu+QHmfrivzktxgS/RThABYE16g0pLugC3AFwg/84/yuOvGVfGyxv1z8J6rlrOS3a
LETxOVYKryNg8y8xfPGF43961IKsQ/+aGDRgWQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Jo4X1DTQTByuQXm8W+X2V/SHKAt5+5N8uNQ87cvzoRW0mpoQ3Hc18CNbiyChL9ee9q7W5nFVEcXi
X9LqrNlNXHoshAD3Lmba3W+7BRExvi1sB4KwDpHEFH0PDEis+J77j8m6WmkxSwWO4EqWKvQ0L3bK
ZwzcAtoNwP0BjWz57maGNayBu5skwCmK94J2YI1M+xVSMLhvaYmJ0sJq4syJ0NB15YqibSTmedEF
c7Nz2deZN34hPbQVtSP+e+B7aTMgHw5NglDx45qlmh+TDf908g/UpTf7hQJECoChz0V9v4mbHbUx
ploW8BTC1EAYYr66OLJ63MW4/vnR3uthbD+hKg==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
JphypdaJfn5Fd6seiEFaA2WjmSvCG6zTkPeLq5P4cDuuULKZOa+k7YI4Ecw+KbBZBfmq5bSKVkEI
620B6rl5AIxSJvga8zFI5hw5duDACTeZkL5YLCt3q5bSGHbVbmGuFqAg/beMkaZuuwCcrjzpXYTk
mDK5jDFydOdJGGEtn2I=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
KZLLWdvM9qGX1E2dLj2e4QqP+S+OlV3OxIun7x0MHsEr7I/1zDetEzNy/awOb3Ha+T+CcZy4sEqi
f3RL92qpeNMRueegzHef7t3um7N6R8pppw439PTJZEeOUpnYKLHGZPzKI6dypQxioQr7X8Y1e75u
0yYDo4S98sRudTjRYeKBVsSKFlBiUNl2AQl7gxtKaXtyTRAXT66pUhd38OwZMa+fdweBBgGm8WWY
TQO2dm4gERK7C1skA5rCsjaoGAvvo/Nk4JN7Uml7R5u+S8+ekpR2o/DXa+3SfLGh2RkTllS+XGcU
HtvChFVF2FvYKUFYDJBnPcgL9kiq1bx9l/gICw==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3136)
`pragma protect data_block
LgWKJIfKsQ3QuzYUrruzC49N0jU+s7xDm1q8FCjVFziwwsiTrdZnP2a8Or6Zbx1HDHGurnC6tJbc
bWofPyaCt6SRAjvjwFxqbsyHwsCNj1MJfk2GWg/qhAlnPTZfcElPgDafMqajVR18n6yI6pnMwwR0
yVeak1MiS+g4Jc1SEAQfB9nrFlZ0R6mqldNIbScw7tikGwTxgqihWYWXC6MeTs52sOELmYUZmS+M
orGIoeAtlwsNIyQFkRd7chvgiKb4TWvZgnElTJmSZ9/wrixez8R+GkeYbteH1LMLE6C0izgTC1U8
VpWjSdS1YWHt3KbArOjJ7FzV+yRsEBMP0KwTkkzM6DVrwSwtED7FsWZApGYe8+M6mRzGVz/PxlmQ
Q8x/BaGazlzBTQsON9oJgy2jV/VSTB0ssY+xLN7xhv2GcP9N/lfrPiP6G2/8M7qCYl1QPhNoe3pW
SClX/IeUvc59t1cBB5Cl+tYdF9Zpq0iO+QTJfO5bxYbsbhYIUbEthJpNZKy6fJJhL3tPoXs6CFrf
dummZkyFnF0AcF18Grt23EPYXgy926AtQbp9Iwts7n1G+xNZDZUeakNa/k/wTuimlE5/YgLIBj+O
PZT52DNRM84o7+OLqI0Q/nDitea3YlkWUjzyBKEsXb4EMDojJXfzGYBj9E/pMzgKjktudMdoMo/e
QNFwEZ3gQgBMBh/fulsRPRBjUIZi1LGFziFwip2fM4gVZSFs50TCP2UR/QKiGyFVQWLtii3doMo7
yvafNuWIv2UdpzNNxzNRl3GPaxXEJ+rTkuroQh4udmujSwpaMzZyPuhDb+GV5Su7K0XHQV7uqA/D
CndlLaUYssJ1QRBiBzHh3vxuBiudT0C3lrAtFhzzgR07khLM1fpAW4SuC12WXxrI/fm2vwC1cYOc
tNwKiz+Fx4dM25Trx6GdUyOoNNe0J/d85KUU9542jv3ZYDjQ/griPUeIiZNkS782q5gZjUzTdot1
FqtV0JX7Bmzv6BVGV0HTuMDijrrSgU7SZGkhlevTTi3GQxxESMM38jrfNJkrCFfWEjiuP7GfSYCt
e6aKvMwBS+35eENnaAiMx/ojQjK9blKV0ZwgIEQfFr4VKFjsul1hNpk+DRRWHe5vbG7XgGPuNJ5z
FEcHkmNt1o//HstxBp4b/k7SqSyzkwNlzpzYWzuqLqNuN60jVEtoWAKAOHOFRYpPtZujfxRFe87O
DKe3g0TqBL7aL+Eg0mU+V4LIUP3QHyc+KHCoT6/9gfXTQceRJIxMs0tGzWd6Mp2UdWJJHbhAU0uE
vjWhsJKXFTqZCR+V4wbuSp+Xa0w04fCSCImT4D7HIvF7WoD8RbeIa6wvaeT55TlqyWdE0TZZpOQr
rsPS7LcAwhMlMyPnBps+Cxy11M3lkJa9Lv75R6uWGmE8ngQCMlp5udxCFi7iQT05cbf2dVEk1+dL
lR12n2ie4rnp43i57ApLzfPUW8BvWcZL+GvXY1Hln29hU9jduW/vwPMLFbFAz/hvUrwqnz/06StZ
rHDSSWDPAwAm3no4sKsmeB4rh7jsIknwspIjQaFvvTpswjhd4NGf6bTCdS4ES8rEJnQrKDcS1RX4
GwRGkkAeVNpBg8Ahc6XyUGKm9pndnmflWlY2OYwnjFlbTazbCVgo3QjAnmGgHMAFFTv7MdZROvZp
9OQO9N0KsRTdQdwTxlXx5UDP3odQp7kAGIwY/kjF1hTMNtVLdc9849Um9vR596DQGC14nyeTBZ7J
b0+TvzCXV90CmiFZYNI51svJgGOtVO0e6w1wNOyLRiWzauOe8gYF1HHn5HYlL6I9KbTzY7pWYVnv
ucOt+2nVqoWlBiIsMGacOiBzgCTvPNomiWs7k94M/OkdZ8l+0wJib2xVSBCkSyOZ94ruFSus5wFj
PjN56KJFbO0stsLb/9L4N99QvTlr7NXoLSX5k9j42TYlfpk+p0F7LDTdQB+nRsQSr/b8vBIjCd/y
nOhgRKAqInSoewWMJybN0FhrSngM+VKm4msupeDwu2JLf+9u4oNkMfYkby8M0K/qJ8aqmYtEIs27
neSQGQZ9u9nas/7adWQOlXyre9wFbR4I/xwBmhuAOEV2SnGPhQZRPeytm3s1jXnw9JZUpt0GpFos
5VJFhbs7Vl8tCdkK+tF7p3omOitZUz/giMPBsKfkzU381pnALz16RDt0ueMbhprTNG6nLefU86jX
DSiAHQtBQmZZAUK2LPcmLceQZiHKzZcTfR4Y7RrJJ8CTaS00szZE73k7/t5fI8dXYT8QjVFwC2uA
tkTqht2zDUmULf6WB+AvTWt8wRhIGP58b66zjfRXHygtfPc357GtuPkwSiKqrfz0ZGrXnN7wx1FP
gCV0ZQTaXyZ7CCZA/A7+qjeyOYFtCBWZHrNDgjj0UREydrRagtfyfCHn9wxfcg+CiSmc1j/ZOQ/H
DAe+tLeA+NANVR3oYC0ZLdfSz8Pn2t1AMi+pceyW4R1Mg91Rj82O7rOQ9CbpYXOSLQDnzxM9azTg
US0l2XDGZSspw89hbKHqCpcFgZqnWeVvpEHDy8RG6XmeV5Rj+AR5Sv16OZNYKbA9V1Lfbx2alCJz
qxYumC34YjuxNICofMBLMOe8GRJclDHvRs9s2GyKhSiGGzPoopnvvAG6Q3oaHr/OazAQkvMKCAKh
IB6KM+dS0Gj7IIcmcupZ2GuixcaIKPCwbmVEO2Sr/+9rjOsVwk2Cl1FNxQT1qFJK8bvzwOUrDOJa
hkYThpIIYu+FDapbghvnn8XRlq6UY/+NDYufdna9yoZAGX+WuLiLNvFa0kPElDFqbS+vsbqvDU+l
A4H3RWLfASkcgioeBEtEXWVOuCop+LI3VgQV9bI+0fIKglmbQ1O8dmy4tIWLpOq5X6Ois6Iu3AOT
QgGYHkx6/YCKVcbPZlaIBuICRQFzrMWEKzDRqzBp11toiB/n2/hSfub4ce800gjTPltMwZz8S4WJ
7B5Kf2dMtawtCBq8b87IRhMFX1ujM4/BmAd4VqrBlBdM8HtpP0cDige0StD/E+cId7MnxX5gjD1J
DFZ/8Vj4Zi7Qt5zDWb1p6d+T5VtYsHYxmvPdfKBppI3LO2T7L5AUnwrwqP4Ox4jSSYxUCBQRMvzl
LUWx+LP0fzt5Ip5U5a4LJPifXMwWZhZoHvP1x7hwLKnKaW5PftGoWqZGT0lMUNO741AwZjbYaWgI
HZJnTNy6HGVOiH9f9+OmL03949kqXOEI8+ojfsQx3S9l4dVVzm/HDUyu+t0khbM/n2IQOQc0u1EZ
vCoWNlaHCIXCk9+OK7buw5HWGsKjTMbc8SuhGyu6htcQnrxvE/UxXBUHTOKkXfvNXpuZVsKtuO9q
G0Eno4T1ZAooRtqpV/tmfvODXBI8UEgpPXRSz2O4SSrAsPoLPyRw7Iw6EAD50YNYxB/YuRpeEtpw
W+DcQCzJI8QGPRzosrxS8s6Qlr1Ak9203F8yCGW/Cq2hgYtR0toHMUEFm5+6y5exiht1oVnKke/1
DSMTIBne+lkY/LI3ou3l0ndQlMXVy9HamIkIq6jpt5e2dQNA1CqfDi5C9HOPi/p3Vhi3SPIG3yGf
wlq26PW99aWsOoYdNKtTIt7hDjI+EXN5cSb7ah9EMHe+fL7DMvEOB5IBpFggpyi3LCrl/mgyvDWk
5x/Sd7tLI94Pp7PpxBvxbuVi8kOMynYVpQ0M/v7VWQawweRmM+LWq+MDSiKaV4v/MyNt767Z/5BF
sEfdQA4B118tk1oLdHGsGC37uPdCj9Lm0fbYTKOZBnCAKBIyvMOPF/cnfIMyh2YZdSmcnEiTsoYC
pUQnj2r+mOBg6hawWwb0zmblzQsJIYRnFbbyO5ZJd9SMO1aVj1epm/PdqnVgXCxrEWPQ6NndChFz
zCGaqIsuGfuet1C2NjFU0vnzsUqCNQ5LQZvD4koNLw41N1gmo9sm5LGAvvyyGTZCb5u3lJm1xVzH
+47OEbVNLuIFpbg7hViv2kuAF6HowLRT004+yt4yZUetaGBWjRLm28Ny1aoaa3LGFDLMCKpCWUW9
LhL1jPZX+F/kdj9GcUf2g6ZDBJ2WP/T3XHOY3/4e62JWNW3YyCRnIpaLJcaGF3DUdtD0Khqlep3b
iZSGp7TE0x6fbu9uq7ywSql3B7FjIErmj2eiDEO1WNPMRtyLrtTUdTYirlr+TWdaBH6tEFoRJugh
MQ==
`pragma protect end_protected
