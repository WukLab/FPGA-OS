module system_mm;
endmodule
