`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
N2VtFTiMai8z1gX50PfTe8a3z8SsUgkYHx76JP+cnNjLvLxm20fasUuicb1freDp3NGoIkA7byNK
sw9UfA8OGA==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
q/U8WY1qLTvBMtob9FMdpIzpqyD7HQss11L6usZnp906ilYvQ5Nwve9EAC/aPJzC8/SLEdRbmiBb
w16em6hGkiuPqxSJkS4yLcZ2OcIf5Mnh0FeAm3vnWfI4d4/9+vV+rIT8KHd+eI3iu+UOI3uwj36c
lLuxc5ahAYpcsrvlF38=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
OVVz+78xq0MLu6oj2NYgt1TP4FMdz9JAj/9f2qes0fKHvHY6X9BuNoh6VmxebCJM6xh4PS4GLckF
PsNhQklL6PvWKWLABjPpudVnEe8Wytzp76GKMrQiba+4Kfvt47kFmZ2OboMote49u76/sROTaZxy
jTkv69Eotg/84ePapg3KXbF5aeCyVAGNc/Td0Wy/yTQk71TQmjJ6I+u3Oi80ePWjKByV8JYgssMz
XEFOPBbol75EaPzMW0MO5OJx6SfoF5CS3ehfBgoE5hEUML6+LuLGwAOuFP0BTay82WpPL/NM1jbh
ASQAutUN3mseW0CLRWOzl5gdkUKvrOOXh+gqrQ==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Kd+R2fKddHvkOx+J0Ftd6otqiiNKMm/dYqyOm7yAhEJ+7gC4MxZMkK9x3JPuPcZPoWci+5x58nAq
SWv+pwdeKOEg/NbKsWw/eC/7jOuGKbMjOqndFqrg7DsGrvlsANr9j/anhcnYps40XLR4CnKHxgmj
WtFmTqptQhrpRr+nPSBKojD5a40k7YyS+eY//KQtXE+85KSzNY2ioBf0Ri2t1Ow3ZW0Grm8chGCX
YhwQ7E2HI+mB5t8liXv+llAyGWQ+Uw5+lQSXYhMbpsH1G4FjWEA8nwx4WAI0eb7D9hfk7mAdGrb7
e4Uwpc7dXcgKjrWcM1VVaf1QlzsPSK1onM7RkQ==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
M2bKnxUvqVqBec94htctXqOokgKr/Tdnvs84o71JhwEvm2qZvAPt9TcKHrc+4FUfRFh5XbRPHCDK
dqxhHlNFinF0P0IWHGcoxSA3hUF9Z5zceWnQ7mpGi8YAc3xmjXqijUU4YcgizntRPfPvN1KJlpr/
4OzUcIWF4TnEXAHTBXrkcihmADagSwkF9goEKRi0PmKckuwmEYE/FFa7H6e0OexliLu5JixJXF3v
yYt7gODgtqppSMDPf+HNuynS1qMRbNPq0xlEaI8b2u1NT+YyFrNGEl5CWAIt81RGstoe1fNBlT63
3ciV3rzTTzPO9bnfmzpFWYwtnHykBxe1EAojTA==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
t9aOeNidwu2MJT7o/0fFm69FSGrd/wUzS1AALx9LmkRdPj6MeRW8xAbUbLHb/n74mMlKAvWdfHY0
9OaPuk9jGqHafqepNr3sJtBGAMxNsZxs5n7o55pYs8mxO8RKIWt5kS0IdUf6ws//IVw98oaT4G0P
gYXOj5oJUe55aRyN5H4=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
XTDm7d4v15wOzeGasVGoNS1jv4qBo1TC3Dc385MNkBeCuaQ9Hc/YMrBjTcfjrIGR2emiHzBOujlL
kLXzxpcOYc7bpxXLSnTUGHgeI67vzVB62cIMa9pP9nl7lKYNfZ602MYugAa/G2EDGFt1xu2Vc3LC
2SMQ6Pv0fqBt0vW84rjolHSfgqAQjz2VgtPAVc2b3DbIkpeSSwwKEMRI1irxnQP8epfIPd3nEbhc
JVEx517X0dlvOuj0r5I+wKIUN3evj0Bn2FJnk0eR+uQ+6Ln9+E7pVWVxe9Cequ9GZzi0LedvunrI
hjqTKMqUyl28rMn0vl4db5aurSNWVxoP3jgDtg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 135968)
`pragma protect data_block
z/vuy4Z/DMK+s7T0lD5A6KQWQt4BfVPhfs4vwsoC7KRdejII/BktgC0uMfumOVwxxvuWmTPjc35V
npHFaQy8JfFf18BaplQovJnnNE3XnO5AvNKrdMJmlW5JQ1I9Fb1T2LcX/assaRjvHG3TpSiFTeaN
iDJ3JY9si3x6OqUKTywShrunHf+Voy3T0xxf+ZryHYQPZvWy7/1hgvTnfT1GwQQvOCrskaMWEmy7
08tF8VaJnn7uT+fMgUPMqCHTqR8dpND3s5Z3aDjlQGRXFZxkExZDfh5CC8gVWhFb+OEs/w4kowOd
N3ftAKExcXIOZtSaY2qDB1mkUNP+IId0oWJMEop4B/1IIrgs/pAnQ9LtbbW+GCZGRY7c2oAeypMs
2EQTZdzI958tmTHyq9LzCJnXEcu8Peu/FhXNqNLsg/oGq5NbNzYpMNuk7CU2Ai0HKLHawrHClMnB
a5Hq5Zvy9xh3siBcfWWTX8jcc2kGqMwjOvjB9+Ca1nwuk6bbHSZwMPceo8ZHr/iZwfqbGS82zCTO
2/7epR1P5cd7KD70k1mlkq6YlxiYxazoZsPPuUBeiIsq4+J/eVmKfUCd2LQWe4j4cyyqVkYVyLQC
hT9ABLCs5F43AQh2W4yL5ZKhgl087Ixf3FaYdCI4Vq6MxNHy/V9EM4AYN/8/RKoSlAtXfVPjDCU8
paWyLxng+fLQJ7Gr3I/yTg+iH3T1apImli/DuubAVU2IItm47lHsQs/SHK+Mf7rXD0CrV8O7Ebeg
Jlszvo/grSFl0dn0bx8Pz+7czXRyOp9s5yaYUAK19CGSA1881mcdcQvCKjNcVqFDLxoD5Km45+MO
q6CPEbbXWU3Wp/qiaw9xveRS53VjUGa/h8ZiSxAAbJGGQkxvQNzG1noYR2mdUCCTfcBZgQYSo2K5
1hMxSHj/NO+vcQ2uv7JNFM0KTPabX0YkNv5HQfWOLCB9htdhxz0UtMq8qNn2JiFNnpm/P0UMXm/d
XBXMxLQGWMrzLWnOBXHntCHKkgFWsOVkz1DCPh1eg7W7/vAmjQ/q2vio3i71uQALbGeHFARTTN3V
CLyPqp/fhdhjFbuuO2k2MMITT3FGsP/7Woiq9FDgUbq0qYhHZbWnyv0xYVOyefDcTdn8dw5Kdo4L
rQp0xkbAwrKfnWQdMZVMCe4JeI94Fm0PVUS/fcyW4uEZQlvYE227IA4OwsUu0GbA19oFL6N3f5YC
t+ueeqdEN6xLuwMk0q5cRKlpLQ97E0+EjlO+cZUdo4eahE8U8xTXeGyNfPdhXjv1WdqWaOF4xtSW
zWoJ/jiJsVfh1dJqyxW2saU9HIwg/DQvn2+dNnoVFK7sp58eTCYAkz3tPee87aIxYdOhVXxHT+9x
fcXbkUWWwl2Quv6fbGPJbrfmCC11I/uCdUaf4E4ovZsoqIJxEa8ZoH41FXfN4H7bbywZ26sS/7fZ
YaG2jzyVHbh/xQ3CiXc78DTNbV3mH60y8vZOrmuHlKjrlETtL36SUJrh5Kgl+8k9cb340stMDlXs
szwX5jgulUKB1yPJb4TAgOZ3N3ZKemTcKtmSG1UAPk0drOKfItBo8j0HL/QVnMsGXMSpGbKGsARe
QJnOOiAbxIO0akou+ASgLUcO2BuHlvqRm+V8pyiMSBnIpuQZ6DTlpdl/tdSkuAQcrKisGV8/2GUP
ziPCSbLVNHaYkl6K7IZ7YzeRmvdK/1riAdJI5Lxrcc91wiCDAZLf0dQF+nTMi78mAXonkrvg4igg
AcmNXdjvaxUArtZgqdESTa3Yy36A4WevuYSs2Y/1f6NV3HWybM88jtLwkQ7kCt37+IOTuqh+VsnY
T027uwmJ5GkF2xyXkO7JPeoMTy4/KvnzS6SwbtXAgf57kah/1f4IQ3cH00+H+7vV4czybWuwuLhb
KyjFe0wcD4acQwNr5bMUe9mhJaOT2nnqBf9atnuBKNpS5MynJWPFXf6s/zTrG8J8v5g/6smkhZm3
HmKWq8x490xfg+QqSccWyRfOluwOltNOflArtlt/6kPqM8jiCMmvDD9rJbJ6qfbAhhK5DoviP7ng
a18Uyt1VDzrGnAGVXu8jA81qwzDcXKNn2EITnkqd/Vy6ljMfIx/3oOSCGQ8FrLglbfj5qD3fELVL
evgQJk3/tJUU0X4oFr0knHT8lhts5hFkU9Y9QHWNbE77Gz4kKytYt/4/vmZZI3GHJYkUTxSSnQmE
A4iVN7vo4R4sKlymLNWisHkSzJjZunCENhihnszda5QdIVvb2OixTNnvnUiYOi37Rrh76QFMarg2
NxNm2b2qUSsLOB0YtgkPP3Tq1DH3PtR/L++kLnAMbCf8EfvjDVsBBxmyyGT+z1W6hL2OnOdejLPX
UL0SD13ZTYPS2B9VjAhJ88Qe0Ofz+8nWiBa+5sJ9dXg1CWaJ6eOJ6EAWMTev4f4YlvzXD9TTEQg/
WYAPi1ppAy7kJDvm4ushvmXHf4O+kAoUUkRcvFk4jPsLJTH6Z2c4BnignF7J36IxPFfdZgwNFA85
5e03MiuezBAxnFQh59eJoCaBTVas6EulGtI1dvENQdKS3omlwr8BHLtVaQrC+WcYGN38nf4+Uen5
T0qCnEKVfMy4mcsltboNlhMGGrJgRQozQUnPMusyIEKZMJ5LwEF+FvoF8a3EQLGXVoEHwokTtjJO
yP2wXQnVM47UG8jPUY9RJJVaH6nOnHDpPPDSnRxevjyitwbqdXYyKQVtoHNpRUoGDmrzO5nQkdq+
qifUu6bzz5Z7r6rlyjUl55vKEx19H4PHMaaFMZanj/gKtMKSxmF78gJxdXcTec6j06mp8g/9lA9/
jdJ53o3xd0hpsXxhtrt7zpiV51AY02qx8kFUoknCnn6GdoQOqNoPBmPFDmWANQmvXu+Du1NeSCaV
5oIzWcWZvVG2WeUQS/ZMIrsZgD+hwOBvQpIOwp655XVQJxIA37BEMNn80D6qJBeuS60QLVCI768a
AXzYU9OHpRMpMCvvMQC5NUKMyl3u6J9ZxpPjymvj1Haim2AXIUXOKr7FociZyyA4+yDXJlSBjX3l
FWoAFYIMkg4iEXD1nJrJbl3NwUz5/Pus0Vu/wTBP8rJrrECpaTybnpUK/fbIXPDiKQDsA09+wGSl
A3QdHzc0+HbEj8/JeYeG6r51c+N1oCTcUjzPnfPKPdi/RynAg0VdCsB6g7Jn45TJ1SOWhJfVOCkJ
tSFRaNXCKcMWtd/+jCd3yg/m61rk+zoEovtKm4BRTH5tE3VensLxYYT3zUeMQQ0WFgo9OSMe+i6/
hK2KUFywPoKkFSmZHFCXrwLXK9gEMdI6dramRNJQ4GjXM0KX6Wxcc/1dgqrYoUZKKK4k+ZCGe/8Y
hWt72VXk+ssaSWJk3h4qEkfIrVwP/G7Pt94s/Yb8N9esC72LDDPscpK7pPHkCZD8zjoeXMlWxlBh
cuCAizK1WDyipV59zeLjJkht0fjnGXKtC8fQTidTNzQtTvysJ8lUbu6tyd4AHsoFPhDO+rAtdWrf
uH7iKRrGq+AzAvbo0PQQvKCGvZxmSEp1hZ7IZJNUCOcZq07vrVeBqnXPliPJcz/bykHPqYkvSiAC
NBI2ggRe7OQk0VrMDbuQR8tJHWT+5unJScWAq9lq6YMpNT1r0+I+uD24BfdJpbMDbc50aUZComQs
h+f910Qs66dVnQEWjXS2i7/N2WCW0OfuCBzuXocPmykg8So2+6jxvlEXuZgjnXKzAbGV7V4HbgFB
DDmgiOb+oP2ANMhklFMVd9IUgrmxpqWt5cwTIIAKZcmpt2TAYMKOW3LHCych/69wtUJsHFlHJJXb
dexyY7gxWG2uUfR54koRqsDDyqHKAulgAyki4LDi04IqqdHJsrAsGpvxGmeyKYFYxAXfoPr7wiV0
EXU2CpXKKl7lI76d927S+wvRPJTk7Buo5QFdm0yijBGlOZR+x1sVW+B5GLNsVfHabhjyqYA373hA
txXzWBczV0NP3HYVKygVWCJvF9k29vM6ar2uqeR38jtHGUxJa7GP3RpG42ih+3RcHbJOw+mi2VAO
s3hJ1Xbv04jN8GjLlGDhQlDbPlzZiplG7nd/WnIw0nERD6TeE3MeOgRq5tbV+P6VRT3j+01/tyY8
NixNS/rIzu+MqZASEWYxa7trda/c9objIVh+RSovMiEgROlu+kOuZkLgmv0ScKDnV3bes2n+0KAp
3yauptVPmfODP7kkCkvyH+c3yVtJvrZzXqGe3kF1P1CySwwt1CY9aVu4e4ZsA5XZ20X06+//y3t8
JkiYkr6wrQDRlDTWedut8knDDzh60oOEaNmjHNlhW7QWdafkjKrN0T11h6RmrPubL/Af5XuVeBT5
u3HDZHoVwk3Aw+c2HeD+OLglNN5R4pIE4EBNvouHTalcFnOr1CnNvQ9/ptyFJcG2dVNmPwwa4xot
McUZQDozlFhJy3zy6gXdgoP+nXBuNG6Y43m/Fz0uslj7acE4Wan5nJoInfIBvU4D6QUUleiaiAAW
DPCPUbGXDQZAt+jOw9c/KUIBHrQv9lm2jvuh3mA+FJxrL8ajox8L8VeRmiIP45f8/O41ILvG8MEO
gzR+Q00qh9nkxLE8YBI3WrJwFx+gnlRIQ77s4QHCjPl1oAuKujrLJfbCh7imQvhPpbXmRmMmh0UI
TkdSjLiXjvSAx/Sq2WrRzscX2JwDLWwMZsx4iezSnDixqXXrPZwnlLs3C/m++25am83H4WBsWt4N
J1tULwTnsQGZkBf/TKhcm3ncH6xSzEN5MKOehqIumOMOlXZbJz2aVoefj6ONbgzNopUg2pb5f07p
sfZ+15Xr3LtE4r9kO0WVC68F3mBt0r1KgJ36tYVQebJUzj3c6sjk4tClwGuZpd8wXCivedm7dET0
ADqfnvMB8qIG1PP2ANVg5ZX6siuGqPnFsn0szcz+n1WH9MxBsT2tarQcznzGX9QzzzsY31hy2qv4
lYrAssYv9KjCb+4sMZQDGLxyfrM4rCnz1hF4hcFLOvGpGapae6R4oMGnfph2jNztpLZAdaLsPPqd
BcclNS/ZD0pCzgKJLeevECoVtOk5zP3IFGdPbEyvUm5IEmf+kFYyi+JB2RSz9iNqtMQRMUtb61gU
QgLC3ftquJLyGSo8pVQH2bqJzeRuxgumw23DSTD45Xzu1vMavxeBIPM+saC1ZJ/h7oPSXLXDNDL3
Lw2U41BjvxYPgV8agMIrH4tvgIwafOPvQzIUNxu44mBbzC3HFDBHlHOFFbOWuTnOs4CZzphuG/cO
FNkJ30MF1ACc/M1Cm43bVlciGupEOqk0g3wR+shh7tfesGGNpJyxDhDeO2Yn5sbuIR4kSwNlBQeb
wzLzTtdTcPOciULqsDUWDfc2M7OwQq8sHRzPgslb8PWVxjQ7q0pAlvunOY7T7otlVYeWekFAmDYk
YV9A0LOi8PEVzLQagst9c5k+vAi5CDtAELSyis9jEiKBG8QW62UdouKnK+tnHj+DWOHW3DwCfpRs
L02erutySaDcKBnfYaRQiNzWSDaj3O6jLoqe5uEwKsMY47r/96fdP1qPqNjBlVRJNjakb0wzt+tN
4Ma+Fzy1mCCPnU+YM9QZO69U2HJSo1sOSHLJabe/Wzc66THSpgmM6+mFeUtHoJaXVXEjz8xHpUi2
n5HK76GVEHx/lBNwW589jPdJU9RXjLtUO1ZMosEzaU3iCU6xiE8T2TWvqy32gzV5QzsVtfdPjnc8
+rmuOqaa/6239aCbx+AGwNA0UksU2/bXcVeAn1qKDoVsUUuzb0kXB8iH+OCzjZfLAHZnpBJyut7C
loFg/gMHdQWuSzJ0X3F4gYrtmjo/t2RdoNCQjEUYtlZbXeIEtXhRBzqFdzv1rsKzbl/kW4QtnUd2
94vf8p1vEOlw7eOdMBfENkHXbQ6zGjoMSC7kfDsyWzTw8+0uurGndsKaqFIV0BOKwQslr2NhLBco
nTmLezsLfIzBnw8+nHh7DVbyUrZOMjr9b7Zrcek4YhLM3jYJUnFTcxbxmCMS0hVXsHvxJrBrxJt5
ORtx+Lr4WL1y9fRYk1sW/FH9TG8gl1zjPLyrJg6Q/DywyK0UT3Z498z/HZMPQrOCHn8oAUINeg9L
nBX8kiZD9aOaLqBHLPe5282if/BlHL3lbpSkMFnk2M3G784gCNShunMQ/+2VyCVYo+qSQ7mzyOOp
m05gitQYFtAdK4rsHtC2j6Y3PANQyZRqlrnqLC3357AJjtw93An61yiAR1rKzoYJm0zlrupX56JT
nOd13AbHcA2JUPyjquo/9an7LQBg/h/3XPafZ7busvbCwtrBuNoGFi+K4q3SGX3P+NCyeciU74oh
ikThRDox+8z/xtsXRlu6/fgYYAJlTdAy8vgH5/U4rGSXRbk15Mx17GmLlkvEQ/sXEKqF09SkOnDM
ZSGMZuWGWfeObBZUwC5BagvjWgaoKqPUKfDB56pIcLOgxzfLYkarWHU8osCscE3qeJ+xZiaYR2aY
HKeewEUI3cg4YE3a31fev8BY3gapjf+QP234OYievD94zxOGcZjtW7rFXgxuGRKnk9EhayPx76AW
zjg9H+4FpL58/24oZvaPixd08UTGir13YrizlcNgdt13bWJGrFGQ8QBf/KBKyWJZ/w6WLkncFHLU
AYnsBolYQFgd/o0CR3nFSP9nt+EebUeKRCJMlR/gNOcv+2Dp/X+aaQ1J8XKYBvvyFWcLWvKiy2bs
zrb6+gmKLRsaG8YqU8gprh/YB5tK/HxINH9Th4/7crpaWBsX/Us5iPoyubJoQ5UNDM2osTMDxxqg
oUrpBpWOKE4qnNK0wfJHQ8Mm0c6lmEDNN7pYRAT5PI2fmvxlLTKa3+vnCY5Qvj6mKxqBzuVuL0WN
jMhVbbxZMqryOkeGci/zmnQkAGp6jB6U+FVc+MnxUbhN1TDLwJ48Fwwrg+NDLxvePA/9QSqy59zc
YXQ4LSFDOKMzQRAGKEv6h7Kc0MRUAiBwgA39N+fYlux/QtvO/yUTdk+DrdIMBDY2vA9w+33/wmr7
9ErHHAR5JZR444E8gsFAqOoJ98kpAQDfTaUTfEA9VTSytqRWB0E2kg9IojW1hn/Mk6+xAAG55UDV
eRiKmWhqRfriJzbvNVon9TXg+gy5qxP7lK73cgipWBDR90THm51KaRiX4OeWFx+SxfgS3aDbmSI7
C50h0jPE7vXmjlFbX0AodpDj4gA05qJetvtmEFpOSEEM98RDDPRlN+DfnCKStl5uRTDghVEzSXGa
rVc6YQ/6H/2NJfOhjFlnxlQGgPR2UVlFkQTM+353WHQZ/6uLwUZKwhji0ZXcDQxvtKKLkJ/Hxlxx
a2bMwh+LQUdUy0mOotHOF7tjKEM1ukSsjdPw/+a/wWliQNshA36/y0JL7RYX5CwNu1a6Vzg/4ul0
xZgtqPODmnW/W5clUZq5ssexwaru39OHy7rtc9a5eqVTSLM94Dg+Jdt8ktmEjmPNnFrFIc3CWD1j
M2x58Cxo0vOpSd+pQIjMkYErJRg7cL4l+FUbEqKaCaP2imz9c49qroZC/AQ4iBVqMgmksOAM92j4
FDs7e4fNzg9lV1fGxUaINxmg7C+En9Qy12O6IczyrUdTkr0S6l1Lky4ucyeP8I8+iZZILt/VMtlf
S6P9Os0RWjOypCggUlt51FyaVySVYm7OPK8FkVOFznS6xUBipPMWq+f0jnVtgfdKV6CxfFLOl1JN
i+UkZ+6AVw8/Sqggb2ZHA6+JiwrielyD2Ch50GlyNm6i/AYOi8cS5MZpPOZktV44mh6vUv+rYLNb
itEWG6XVZLi8Q1YmEPuOvc4gcc0Drr1UWgtyQ9G5Lt8eUVJNQWEfMNJ2mgd6a4GFkK6rPcJ+8IFp
CxZkb8XUS4GkMYO0YJ3ljgLoqBmliNy//OPd48nBFDmo/IMnYBxNCDT1oQkR9xXXhMd/6/7Shzhg
eIiBLwr2JwTpQ6nDmlgVbCYLiTVJpLqs5UfoLgzW9hlMNERspntYJZhLalt+woFJuteznLlnv5og
y4PsKkWc+tLXXaIzOY3O1LnSiPeuUtctCI/QLilRV0xAAUwY53h6MJhxMhIiq7Licb1LpLvdEdxQ
VAx6DiiNVqRLWQYfn9a8ylZkVk1gFm+ULzyOPlW8c2rIM3ZrNZy54Y/HgtlvLq7uXEx1K1O5CY6X
JIDmYRM0uMbK1jeL/GYRlmEf2tBn8CvT7miurNz5dp8gJm0Nn9k0qAGrCAtB6Rib5ko0U6HHj70F
f9su5J7YxgxGPzomFtKJy4DU49Kg5ZKdmdCdfZRt5WKjaqeTn3Mvf3CIIggzIZh/B5WAe+GriAb6
LuCiuKvvd8L8TRCllHGgilp+ZuMXgm9d3pEqOngtVFtb30mWK18psjzHMd++vEwh579STKdsG6hp
1Mk/eUI73UHZ8KB3j4+5IksoY1gfAIqahrx5ZSI/i6GrFcuXKsNsRuXYeTTugvzRhYiP7XZzcoVe
ILzh31j7Ga7OkpPzlwIUPDfpmbJcR1uSnY8ZMGO45fSSJscWBwMeX0md2w8wGhjIlMJQ6unR0w18
slr7S60XbCCjJE7Ckz2ahWNMM6lJjcqk87ZqTX+1OVtJnw0mGTIj7vOf6oGY+Cu9tC1rlmUCfpK1
zVN9l1/FWOhSdXnlsUpTL+7U+McQO3UWeBdKY+/q1ZphG71zIUUX7unELj5Ftklhan6zA/HEPmVj
d0D0pmGrsa8ar8z7D4aJgyqIskd+RKFSnV8HHpJHhR91juvXHq0xtk2SYVsl4R8NvKLKL+dwjxYA
wiHDZvE4205f9ns4zGgYnpJT0YgMraMgHHS/DD5SZypMTOONedOlc1K2ThMRFSfkcfhKNXl7SRlM
qrrhhBXfwl1NJYtjFwA63XZPv0ppbSzMh7GHht9WGCxcbhlC7p5bggIcOiaA6UtgTIZLe83nrfZS
vkdOSJnZUvsxw4UUY2X2pcJ8WYZV47j8q0Y4lY+4mazNp9cEGz3L0AEte11IYih4WFaKQimznGx+
FQP4yhXxk3Z2HRC6QfKtlYRiDBkSseX1d2s2S89rfWmRkM8mrCioDGhM9OSkfy/+Lll0zLmB2DEW
21wVRj6Pp2oESlQe200AaR1MaWrb+9gZDetpuUd5C6qfs3Jza1xOqiGjGG/d38JJFU2+NwqE3M3s
Inr3v/Bg/9aLkpQPD7r/IU8Sn0K7QbYRoV94h74vDuGn09sNJVXeDXDW60p75diamPXg2NXnPmjS
Kbl0XmS76C8U70vVt4H/qd83GeYEe+L8otPHXtttWOWg1cbhsfIJsYus8U1H7sCOI+UeFTxn4QER
ixocpJEsFTteUDIotMkxPo2uSnabmpbDtCJEBe5l9b4EM60zbDOkuhnN2C4vJptSF5YcKTJ/aTd2
c9XDHpbWnem/l/KDiiuclkDnXj8Tf682mvKQ3YcaaBx7O1Pljw31E0mbZn0bZBIaa47/8zzteql8
SrRVZh8jt562oYYvZePcV6t6SBT/lulAkyerf+6OtT37qNxtgoG+VccLjGEFDkdkMuAiUiEbBS9V
xNGIOzaCiuCmgJ+CxrOGg3mqhMWF65deYeRCfJMcgJttDPmNzvQLBmwg/w4cmUSR44904N88sDCj
x9Y7zwLEhx0doJntDFXoIoRSA7V1AhTdujjsvIwFUOtl6ViAQeOCI1frS5IgUYjVnZm8hC6cGEvB
YcL4FsKm3Ai9VeI8jH0R/urkPIy8fluYc6YENRdnEIztW/kYdLr82Bw8IKW4GRo16F0c2jeyPFlt
HLsZhN6pK2GDN8r+nOW3cIbW7q3MRYOFWeuW9Slki5+t7OOmihwLrMlmPHfo+9nS5Bde/fryHVCv
1AWzSswSghq4FoJWL9abam6VzHiw4oc3YIzL2rwN4SQQYfybMbpMQb+9bd1KHvAERiWoD5vv5Yfh
SS9Hl2Ea07tU3KoTvLy6M6OciOiRM/a/y43kgjpC29o2kwiqxJR/qIxPSPZ/KIRzTP0lYqRH1ZQu
I47Koq6NcSP9CS8xQWyYlQLi598o10BElwWIdTiFvrkICkGO4Dky/9WCAb5G/OYWk86VtYva5t0E
TYEXPX6A0ZbuVSadFetp3XH208saPUl6RJPHtELnR5BKvOPnh2PocCFJD8UyEZMRHCcxv79Bwbyw
NrpNCzFVeuy+IW1RPq3B+/Ow9+yBn2LG2h/Oy9gbPrfUk8Y+K3BGm1rNB3Pj1hMuMlNn4KVYRPnk
7I39wp0jO09Dkoj9qYaKnQm3aaT8i8rdNCZVT6UcKev4FUtPyTknHmM9vWguP37GxVlv1QYeG0NB
Mex7CNyuL/XrclFc8lHZx/zlN3JY+vOhgLZj++5MlJabJ5ZCaKWTYwXhiHirQWX/pREXgzJk3B3K
WDYV5I/n+/UBZkWolz5eErVzfGuAcbCROBBjh2bBtX33MVzkPcGawZ4YDMH4aEFWxhpORO/+SrSO
eSfWwG/K3v/GrUEQoqVFEhPkhbaaHldstBWKJcWNApZw32nSuFWr1/5rAUppLzy1AfhT9eXnktPS
naBCHGulqmMGodSZ7E0u4cGkTUW/DUQ/Z/24FC91h4FIU8tTGxlpkT21q6+tQfaAMei41wOxpE61
zuy6vlPW3tI4Ewb3vmCkAykh6S9EgYu9CvkSmM1jHKgGBjGjG+usCsfNYJ/df96o8vzq1aZ4AHO3
WYpFHc+RiqMaOAWYdWjMhAINVUgy1ttQKTyDkylfx08HtfGKZjjXKJPrKwveweGm7Q5dS8K3E+eR
T1nx8JrB7XhPaPcdQTpRfTHTfY8yTwZ1ml7H5cAaLUltCVGhQp1TT4HqRqt+5INzkn1SIqMDst+c
b5viFz0CcTTAM4cHsVrHbcxdyVRB1iiVze13h8r0FbA4OYsuxLhy/5deG3BJNt4mVsOIPSWTv9U3
8DJLrYKGERdOZ2IVLWKVglI5yYU1vGtEy9Jl6WBGRoQBgU5+qHFLRz455X+SK8+IOkkDROOnB23W
blZYMEM7Dm+qcuvU2b3ajYeDTmK6FAmNcgRk3rEp6TTud27spDjWl3dE20xBBap0koa5hzxQ2Eec
+o2RT56bHdwJgz4ePwQiEcoU++EQAesxDiswf1m8n8M7BFmzLYobps/ZnDdZqXf+/Y3kG9yppT6A
qNkMMkUHAPSZ/ohEImzy41G8umrUvOJGqymLxe+YfGhUyx0CgP5bOU9uhGjPkv3JKVzHk1j3jido
GOx1bCoSkA11Qpx45uyGGCSteTwZ+ZCF7UrPFeBMWwrKyxupo2leQThFzJp2eButtXY/8HowmBl/
hBjQz7nEtZaLYyaDzFgxX20oIctZh48oumPaQ/Mhe/NegconOOpn/Oh6zA0cBYWmlPjCLQnhEoek
t7M5/f/MiKcVo8J00VWmnCoicz103VSOLMBRAXAJE0tlk+TY91n3k/O03RGN+I2Nkujh06KVeIMo
a9rDCI9/+4iw7hckliaP23p9MibXSsNsZqvq9fxJzFUyl86eVLeH4n7ADfYlMU5FzG2yV/BA1D31
/e6fHqKCoj8ewJw83Dg/dq6FAp+Qg+dNAItqduX6P+oiRtUP4xbVwf9lNvXnyryahNcqZZzGDqb2
pIklpE+6OOxoTAWaJA9t3/Rm4J1wNU9xD5YEYgPIfSeZcs8DZB8/SeADcPHlpKfkeC/yhIlFplgO
6HB7I1J0Ih1PDjqZWhIEERZylC4ovnxuzxXMnzOOBGXLySylso6WsD8Qr5rUeEYg+yUehf/rODzz
C7MM1wg0TdszfKGKs/1qZ+Tc8D0It6AilPlsVz9vRGe7YuZMda0g55yZIcplMt6Jo5WX4AWUqpU7
dq67ksGRVwI9idsV21S4cUKwn3kksF83vhdLD0hzqLICj6VPPNlllCbQWfrHfBlH310Abh6yIn09
fG0MnS0haKrqOoOGxG1EYxeE/UF6OXK1FFSBahOvqgiDidWoYTanuMKVsKOe9/dtLjPiHSSlmQ2m
eu2x8iB5mktE88gN5g286daY1e+YOHArzfxZjg26U0g8Lz20R5yuBILjWicomjP9PjT2Oq2JVB8+
vdr8nhGLcUGJwsMvBTfSY4CdjpLuwamH+Q09gTgeAp0sfUbnMAkULXK9Huokwp+iqOohsyrZQpxj
zDX+kX+La4mcg1/0wKA3LB9z6LTwpGiYH5lx7ySEeorjbOiOAXioDyO43ZLXTtCxLjkixWQeOeqb
MYftKwnDg8W4fIEDSFsCAoKrNVrncBPkTJNZEq3P/n4+Ue68Ege8mR3btmYQ1wgUIhStkAlyyVmv
RkdWn5jqPZCItzRplGZJXPRmHuOs240pfvPtLDBLeG8mECMWcrK0iUVAyIRM8C9UpK4DB7BzgFnz
745NeTZD4po6xCB9q2fcWjrnik5d/PFYmru4/rCbiLK8DhHmXoZt5AT2VT+eaYN3dDaJiAJ6ULyp
tCDNFJgT/dykpQz5R2TyzTqv70tbhvOon1Joexs3umXz+3/R9XAybO/MN4R3vFtJJxr+v1Lo8RHY
qCgo10AUNTbhv4wZRVVxwBWbhgAgwsDioiHGrHN6Qr2ZUm8YjJhydcSNX3pO2T+OiNdiO6jRvyuP
5Tpj61HpEEjpIZNDDDAgLcPkN3fesv2t+qP4zjnbc6ZsyJCslKY7WPc2eHO8SVmeUO+LHTa/2imK
cThJcHEKzTT/r1otzSAfMp6m3Y/FN3TSfhpt8LLQ5wdh0LPyHadyQlqaeeLkeaBJ46VsAj8loLvi
ozbt9/KKfmqhX/jd7EHrDRR413Z//+z0EOnSGcCdY6PAl6TvYWhnAPxi5ILNyaBVoKiBxaMjdiAT
GhdHXkXt3ycIAKNs5NZJE7M6bmhWyujchwnpGuoYAZ6xMbbJr2LMnr0/px8id/bFRkDwqudOyb0q
Mdm7+laLzu+pOiAa4rpmrElGX2svQxPvzEngJnPQ6aKuoAyv/P7yyBLLrxZbcYOIsAAkT7Dr/4Z+
tBz333hdj3JBNMM/V45coIDAklNVxa3c2U/T6PVtvcyNFX6d3rOUwSSx8BxE7IDblHhUoZY5IMkS
pPpr0585o9nxFk7bc/G3C8etsEHWBUtsrIit8henX/l0XGWwDE/6IvuS7uTDDGt9JXRm1Lva8zGa
ZEngJb0YTmP/XwDtoLwgsSPm0ZEScu60yiELuOydRNLW4WDTM06W08baXaX2Q+Aogx1plsKsnCyB
rw18Zxz20CQiRMJ3EVe3BnTIGL5qII87fg58Y4H6PtMBVf2Obp2HLSnQWZfN/6YcIZPuZKrbA0gR
eCYXAzRPKNmnFrLNUmpHQvbdHnw2L/dXl9IShm3gVP8xiPDlqwlqQQI7n7wmZJlQZxkl/sXYbLxe
cyUXwA/txdSGOZdnr8xNf39wBaIYsKckgtnZ06+BDnGoWhVwHnBI/rcIdnUWnaobpiQDoQEohT13
AFwOu4wcFC3+hDe1N522HxEgq6nauWWlB7j/ApXeiGP2Pwpt9kcadBsDXy/CWCBY+LPOFkfT2UCY
jCnIyW9YPgmFeuckDLQnzIw05qVPVS7P07sZz8f/DLA5Li6mqeDg3s+GrkQi47i6e+cAh+MCUYyC
8be7lqnEmO7BNa0Dd6k2qUoAVBLADd9coEdO+A4oGa1Wm+f/FgBpmnDkfFaET1bdcONcd1vJlN+H
Dgwm8D02+NFtj6wH6Yqg5gwqBeAFAZNN5jTK0C96/eTKiBr3pHd32xzmGrTPS+s53tVP4HqiWR4j
dzZ5Ap362hI54xT+HeLfuLLSsQBsLGSz6n57JHoh12nyD+p/uZGdg679PR2JntGQMsMJhA6FKB3M
hW26N7GbQeHWqSzxCV5fgeIEfpN8Eup8p3QMsb0xVddeUyFJybXfOPXhO4ClfFD6hy38wsOe2vA7
AFAnGUdAbtp/j4b2yycaGbrkEroZJNKC+EPhgIns/u1K8HD5LHJEo8cXpOJr2YeAIYDbzwpl68Hn
X8B5+HZpxe3ZCV8wjLv9l+rHRvmTFVAJX8UqRxcr8NzB91fbrIZyBhfqBBZm4b4JHEQfgHhKhFIi
gmSKyMqoJWLLfypZIilC93UYNa4P/PqRaTT1dnRaLM1wxt89pa5x+yZXGQR7i/sgRWbipjyvSZb5
xZ6t0G7D8oRPD02NiSYCbUUVCiK/VS1ssMTUPPxz1ZCpzSSxwD/+4195VKxuwoSwAeOoCF+Wopzh
RTzW1MxdTuxrQqSyaEbphMFSOh5D5HnE5u6pGpRYMEtUAN2XtGB2MtJT4oLdlc1zdLjipxavRrzf
kC2PrFJj7SYGRy7a6FUeM3DHeW6SF5ApR3T6GILaufXuHq/xkUA2wZn3v4ivrxjnCaDPlasLiDCN
p40Ks7zr6H4qjZpkgFAk1JtayW5xgp4lYBdLTghVbXPA/EPWjJ4c3QssBbihVAGGVDId+kw4VRZW
zc/d/c4SktqpXYKk9FRKlatTFGAky6PQiGeLNywvR+PKELZwg6Ud29bDAEv1wMd+pdwgLqygwj54
hrwcGK9bDZLoDENAoc0NZOaWyLkL9yXgVF+hBSI6GP4gwl1pPjmZCrj8okUzIuxzFXBIk3gg/oE9
lPurmDy1VgkoMn+ADJbUk7b80P6m3pa1lchC8hfK7IMIpLKrZ1CQwuMiVGyXa1JzxBYUztL4DtpD
9mRGWivtmwptovVospxMAWym5RB17o8TbR+Un3D6UgthbLC0xkuD8mhXlj5AwMlDX0nixr9vpXuF
jI3rIqbnsAX9BiFsKsXS7iquWn+vKrisNMluEhVgLDsSQM2ROvJG32OtaOiw5MFRK4g3yQcLUMRA
ZXIlqvUxJm5RcblHin6m/majWdMoe87n7zIHpxdRnoTgfW1naJ0uCP6VrzxLiBbw4S/2F4KVjQw+
6ZH+++qJuAZRYkv81Fse7IqvSJLjiLIE9gaBkVgaFxJpKr9HItACR6Nlu55bflEWOSnmbVkyn4e0
Yvmce1D0GlCWkyQhGs+V8WZPEsOJ+Os4YGE8vOjNjiOe0sy/9RE8vipH7CV6fxKdGfG2C6lWMZOR
cr64zVj8EIv9b22m9R9WrXyldIKWkOGoN+kcJPNL9Q8nKMGWdqEvPCFzu/swbz7IWHMhvgE3hUzv
+4C9H5ZJWRnMpLP7OsWCIhH8O+5/tZzgrACwKdYrSY8NQCxRoyTs9BU/Jm044fMIWF6mnEgZ1CVA
SZUi8Q2lJEK+43yydja4KaSzXEuPEGHTB7jsPBD4bzbQBNiYcCY+zOS6Qicfq71MWcNe5w1gYMVL
uvNBQ4vPQnD/UsyEGuEMcwhgWVa6k3ZGM8mT2FBA64jW6fChJPb8Vsso5aDQzL9Noc1b8aqJx8xU
y8UhPrEPVHwro1GITuxbkvS1WpD7NV1qbKCm7MTtwhakp2ndBA10bJ07LKsGDafQZYREftggMYZy
4HB4uEl/lIUkYJTof7MOPmsAlBNu9igu+IznYBqWpm86dhZbjuKf4Pg2K+BbZsoZymrHJW+xDScx
OEeHPudDKVO64I89r7G7a3G1I5m2UwDuzHUssNLdvyjdjk8jsyoP6wkdpH3uDJkf4vmzACNZzy9I
lpl3Ny4PSoT7z1mOrwnQF8LhW3S6FoDx/Jz0z88v0tD6WyIcwH3EVEL+rp8+7p9t/LhDC3hsS8eC
gGTTT/qxA1m6ke7psPpTsF2ZeY/TGggU6QAuHVy06ltdgknJjsPqPThqXU4UyXupV7u242dQNVXL
FT06vkrXz0wBTfcCuqKVLhbwN09woBlied7iB11NZg7bby8Ii+O6VbELs7NnBOm80+gWXPZj+qQj
pczwhBS/vtEhTX+2rCAwRSU/u/QyicwiJEKw+F+ZwwazbFCnReHvxAsRm5GQt/FfdVgzQsKpSNzb
wC7s/76kaTa9oaGE+YaoyDlo7/r4nfaOZbN7MGAU63WX7mjGFNyyarw8FskCj+2V3hV1NJ/8U4ap
QE0xdbpUqxIOyeUWu5+8kGAa+9oMVKUnHJC0Ra70sh/GG4I42VeOmBodK99XwsUh3mGYxAtOSKhy
xs1kKnXTzWY0k51Eope+wzxsHFtk8G3L8K/JaZr/VrQQzb+5kVrJIHLuiK6yDP5Jc2QNnX0G4Jxn
kODnkHPhBuP4AxES9ZVRKXa/FG9uiscsq5PK5f894PmJbdtZxkU3E6UPRFlkLro+cVk0O9Oc1mq1
oKzQDtLE7VXGPaDOYf+NJVmKHOMYxk0kvRa3qUiAZ8EaXz+lmUNRo2TDMaPZUjFWJupJ2MzqT8kU
S7jkey4Um0Eqc0v2ukgHZrLjWEY0Po5socKUdSrBYPK/HCe+lkAefi5YEuq6WRhXfjrFBpsufPKs
PRurqZU3C0MKqJTMNhwbet4uWZqvmA3MJpVpeaZjRYvDK3WMrx0PXGEnAR9MPcaC7V30Z7Gabs9m
MPyGpRj2ijqhevIPy7a5vaWPLvTYcD0YEVMosEdhNrlI1/E7OzvQuzxotvwmjxOdhlS6HOGizfp7
JH0SAMQZEkQlZ45AI4+nSYAT9yUzs+DWK72n00RUYgLMc+z0UNDjzJ9Rc5V/kHoPzAxKLKcV7r7t
ysG2oM+NZbCANZCdNHNZibjNC9I5qwAVVMl1g6FQ+hKQYZjYz78z6DfzDPY5vGPrqoRIf4yUfY+b
KeHqTWupUcLFseDVQ3qfMujms34wj/H+heAQaXoMf1NNndwwjcdMhQd6cn8SBZJ/uZmiRubPfJF1
jTXxh5TBRr6fI6ewJyOTxyp7cSC5nKkPrxhT/G+/upZD5uD6FPF/yatqx+liyoR4ahQzRWT3+bPA
dFJmtN1JtxoY0P1DBcMs71KDNkb9P8zw5I9HU+IHZ6EOG11brvOcuV9+tx+ikCiPv33zq1dJ6sdk
AKh8uuYZFPw98rkTwy0KhG1uIPVoobGXsZwWZXEpsfuyCVeW6TCntDFvNrOd82gRT/XGZIMtaylq
mKN8ds2APla+yomOcWMqtoOXxd3NFJSE9msoU7FIMRDUAhamVBabohkFvTzaroMlGLQqtr3ndKRV
qw/SnaBKyWoLYBLGOZVpEqdo2TzPENAvJ375Hv3qejpTt9j+QN51f6b2VVebwxHzluPrwdTRvJI+
+NNsG+1SJRRQN05iKt4SNix8fUK6HDW0h7zuLzvKY8BruhFzsT6vQJj7sJx6ZfqckHDteK6CVdZc
se7nv69s66oWDWGQ0EDEnLWobFF0Zw8oFTs0LNNP9LPKw2eMfVJ2uJLzHlt/iA5r2U+kLXE0VT+5
iYPPE/REERacIHAe9uYukRXtUTgJ40NTqNJiluZc9yW6LgcRDozIGfhQbnigfNcApNhuZU2NSMUg
v23r1OLhUloXhKM0oFWW8EHgWpkbVefA8xTEzSKxrbDBnV2b4pdtwFhZQcJ0WfXQBLjKu35tbYgR
fiBytd8jCJXfBghlTdVyGMol+HIAV97I7AjVy8Z6YnfQR5DS4KfBriDW2ySLCkneepkrmxscgC2n
q8S/hgk+Poq2QWMhywKnfpRf/L8r4JzYB7BmV+a+G9xyCaDl7w7jQO+uPNtPUd5RHXQxrGyfiUMo
qr8EGLolBnBYkLI4YOZdWrxzT+zJFxG3Oc1xrqkmlAHarQvUpDtaWb+/u3phyHSQkaYS56wNKc6x
WXfYpuelqAr0M+7pWn2Pkp3WANYyKu49lN8YRiCx2MBg9VZeQAH1LHk9zeDu+LGE3M4iGD5nO5dD
0Uc0YTi66He1RFDdWEf7kEOW4N2l0EH0Ju1yk19+gNO2mRGm5kvH/4vsHBd7piBxAUdhhWXXOJbb
GfVojqwr7NGDvBaKUkcPqrHeSodw6+0AYWdsWMG5xuvIwOHTeAUoJ2bAPfdstlLj3g+qM5VoxJoI
UPvfXCAZPW0y5cwzyUcUUOHuz929gYVditVgriYOr3quvOeyQSmB/LvmzLIDUX7jXK8Astnb27jM
k0uwfCccSnfIw+99VBaNPYRWVOjkrlmmNIgUdFZA/7j/LhgUhxXnOX0721QygAw2sezpIeE5heq2
SeVVE/RGRK/wEqm59UQh+FcGlvbS+ZXxc4GNwgsRgzX+vQGzmPPFYpXTCkNdDUx9YcM6AgxgVY8C
Bq+vsTcTbxcMlQEfT6HFbfhohJKpc467fEZhK2lqSBR+gXVfxZv6+r1E6NCajmaJCKHUYUHcCk6H
/n/nrdWdVnzQ9cWUQSgcNIIfjSK8j2UrVGq2hWqlF7kP4HWTNVlGPqzWCPhPEjvMkYMte1aTY2Am
w9Nzsqr/0M/mXt7F2z6TPYpzTIx75FdDUsLF2IsUw8qB0G2SIrFtIag+Ud2THXqe9ldccsOmsdog
fYtPIrN7EljabLB+tCQhmdRL26CVeq/rbYx3WFoDQyg4Cv894sO7Gd02vMU6TTjToB8c61lmm61f
W/eGOucvKzdNwLCE4GCmI7lL1LFHeG6gblbKmRL+Ll33b6zhm6Rz/R+E5ZfhIFHplaf17vDDgMiB
VvoXC7V1+/qP+3SEKnzzHnSlFmyK16JlHR2rRE50c3bQMpj7QVS84/jRs0eFzeN6NUi258SW9f5E
/8fFLV/9XiHzkKN48wKyghh9N2JJ7wJPna5UmBFXFC5WC4A8GP2yMxEYoevtmY9kvxwY2cvUsYes
ywWk+jR0kjQdChKb5HQ9j1HApFWJNfntGZw5wzI9iMAw4pxMJMLYu28rCE2dlr3ikovQX9KFdwi6
l6JwfdLM8wvQ/DeB8mP7QNcjgNdDe3ZW578m5XWMuj6mkKHePYU4XVEhIbwUr9WwCL0TlWl2zKGb
5r0FSVy1uO3Xk9f3QoAy5fWdEPWZc4y7PIu7pwCFXcFCy8h/tv77rOiz4QK9sn+gcJTru1bIkwT7
PtgyVyQMWssVjbG+Ih0uPB5f/4P89v5WqwkKCyQn3Pe8VfmMVPkKS9qKo+1vg58rg3zEC9vegXSX
a7nBb/8vxT80RehAIvn2wl83B8m4xl9Lxhc3XFiNCvS62TcGlEsm9eVpKeMDd11fclRxu3SQzsh5
WfDmr3I5zdnP1bP/+qSBtLUPfqZYRMkqFp//lCgpBRqVjxt8OBaoePpYrE923p4GDt2UtifBo53U
BVH4Go/oHnV5ipp5S+AUzW0ogG8XLPCAA6DG7AH49c7p8/kAtgkG5DydbUGSPMabFeLxzWVvkoqH
k5UD69FCfUqPTpkBJspWQo4GcLG2ZUi1OwE964zkYZZgYJ7mQweWo61f/ZUDw9PGIIK/l64HsDP8
ZSGhDOvOwHk8MS8Szt7vOqn4EKw40cu3HEw5QjVjscLvthYcSP/u2uN/H7/yuN/1oHEbkjsT12MM
nv9ZWA6p4SHzO8oCBG51HqCloWMFfkp1utTAhn8/XRMPnRJBFYe5lZF0um1KEDitphIUhSbCGT87
wQsyuMrtewa2N2iRimtly2UeDrU1aZRsC5rlpeGEQusv+nx3ISDpGOc79NjQYnR8qtqjtgInfXSn
EBx+ebEDNZNVK7ln47BJrxEFTQUP3ak5Zt9U7PN4MjJJnrB8Og6O9/UTYGs4brgrqkqU5jCQvr/m
kxSmYukPItesHVppMBG6Pug6cZ+AB8ySp2D2imPZcs1/H0PA0OiDEfh9C1zjMZlmhjMj2Y1Slld6
xR2pJxI/lMwflskupAZK1ki3PIF+JHfTY64kAK12RJikUTE1tuCfNsL4wmBUfL5AvaOLRXfiF+Au
c/+QgHw6mHal90tO9KmaMgP7gcBRB/+LhdRhUipq8eejlBvfH+xQon9XqVgpp7WIJ32JMZowVIPa
cNlcIETfQUMlcMPt9LNq/raKKAAQeSv8ldehmL9EA8bgjs0VE2h2UCEE+Gk4gGflnPzJA5PdDxEG
KEoqUVBKLJEiiD1lm9V3CndvOmyfyL+zf58lG2yLysSYZphQAxQZFoS6zgrnGFmuDF3KXeTZ+QgP
dbzwEYD1DT3X8TF2ZyhhnPDs7RWM9aqbjuugPb0i+0ykEqaTZzov5qTG+GSATaViNQOApfcrDo5Q
nQt/uQsxu0G2OmL+v+24hxWXEfj0VnbVJaJA6eCZ3KHHf2NEAc5fWuBO2btGAy1/gttPHLokCZ5e
PkfBQ986kG+RyA+jyRgduNKJ5Shb96IexJItKWU5NxJhpxeD73gN0KVkVLe5n0qvEUFkif12rU5h
kXVOrU3jBXl10UIzCz+eu2ckhQ04xobzvt1hZ93goubzHF8UuDqzpZuQs4pCqsgocdx9Xr+vwW7X
0miAxkbIcyi6Wi4QPd/Bro36wUrP9nAt7KrkJFC9DuGhcpfx+bTFrfXnm/TIyMHxMBWoEEvCiEa9
4c3OR0UwKoTEaYgIEDtDZGl7VBvaaJmaFhGRtYM+Nxcnb916SqiCRpql1JZrZMdb3NZsy0cpOhVB
p48kCEmHYisnjtP/rUc4DnkkASrLSeXRrMp4kM2AHOn31Gh+FfP9pX0hNm7+PNMRo+SDe7sg/IiK
s2XGST8SGw8YDJ0FhC8wj0ChlevRW3AFQ3/VBpzFphTZ4XLL6IGLEQ3G1VaGOY/Z4X/tBcl7SXcV
E6ngnxrQKjC//S+3Pzy2BcttKUpUuzKafkJhd0HTCY4T40Qe2LS9B3CLC9b9CzmDXhqUkfI6CzA1
hERj+eHHw9spnHBLcrm14XM2ZQb2ZL8ihvStWLrKNCBklC/A/haAzYhWQyEBbkOdqkhOBtPl/AXN
k1eqOBekcimMOQ/IEZKZQUd58kFy3AvE3D8BuZbPlCN+lV4EUHTEeDxSOT3+MSwRy85I6J1Cj1WR
WgvwsbsbA61qnemvH5gkSpr+9E9y1n8XzhBrjdhBJx9/I44I4K4HXC2iIBSnO1tw3DV8wbhWnuaO
eh5gCdPSIvRAn3gjsw8nKCud076kD3Axu1B0+/O7nqkrBHIf4VthCin7je0Fr1+8n8Gy5JnEyqLW
y4PodGhw3pPz7J2emTDMO2MV3j/kLaJOiqTGYJqUuUWKoWI7qH9CwNLFl6fQNwe/h6FJFZvahP8R
fqZbzviWvpGXSVXS/EOF8v5LCZn6TqnPB4JMAEXKbw9pr+U5VYWTruazE4NsTnxw+GKPA95RxP0O
nLl08yBXvpk7O9K7Dfcbe+hGCIlOM9KEvCdaq1MwHDAReuVsu48PSw2y+9htMGFExwKN5bvHLIFo
lOjV8p5eTdTyIFo7eSvWfHMCryeI750M5IyLjQhAOh6+R/jKUTqGDrphHr4GcwOw/pvcrnYfkEFW
wD1XsLl6t/JctobtQ8UopZoTUkTeXRHYf138yYfEzSCfbHXsTELj/vlGgNN5w0m1KDrw+YXIgOwP
XQeToq1aiiPn0mL6RefKs+tkacnsLDrnvhWkrOAdgd83bIWxyZxlM7444IyUTU5pxrYowpyE1FPn
8mGgL0Z2c9l6gpdnyEMInSyxT0aiYvQ1BXaw6gGt+hiY5We29QzpkSQsFrp8lTFJ0ZXC9HL6pk+h
HXKZ4+P1BNv0YCG+2ai8I5DG287elnSCOlMRKWad3S8yRD7wVPkPUdLtU1ydmkZP18Idv9MnfKpB
7+5uTofJeEfoOboVrZBvs3BIIBq+Mizl7499SXgFMifuE3hi612XfC4WdfbZguUwospByldamLQG
RGQSQ8rQcKgr5B3mNuscevvi73PXQ55gLlHwxilKwowh7V7AwRuP8biFub6WaZ8u1yCQ08M7xD9q
F5YXXPE0C2P4o97B0G/3eWHmLG5IdsAbY17mQzwTmOzfcnPrpUEMOCTC1SXxPdxbcFHH9qcX53vv
dwsxfNbS2A0WKYKl8zvM630zhcqi39C2/SMx5Hn9hePPUpPPj69mQSkHJfRklVOgOK1Ho16YAI6+
0m2rKdCkMkkRnkg3tejucdiaz4RgokoSdNgAQMZHe0DBbIpAcmQR6wiq9yvhRyZFSq1sqMqlSCkN
Nq/0XWBjEniSDf/TZiXACblrxWBuHGG4E4JPawMO3Q4xfNCttghv3Za+2WQU3QTIGzv1A4EpXjSc
KHJ+YaaP/wuw4aoZ/vAB3XIEOkwQWh2Fpdd7lyWvyvhDczNYuTlCnur1js96018nunvUnoNFgeoH
I+gota4cEhQQTY1uRMQRjThSpxRpQR2/skGw/174w0ytZFCY+W70Zq4l8V8V8Apo6BdEuH86fcdD
I0GEO+VYSE/3IsAyf+oTYsyUUiADZ66Sa+MxWf3xSC7y3BLFz39RxOdQTiuj4xkpsvo+C/0ceOJU
CpIIvhkGCq4BCcfd9MN2QYFItzJfcJF5K0JRktKYpt9IbwUnjnWNDzZfhxkY7eejFGN0ejGJYzh9
A8++MFwnFPf/O4w6NppFcvfK6D2MpD5k4nTK4sF+WKON3dyTpzrW/ASkTAk11rOCpIlVMagrsfS5
nuuKMpcbLy4cxM6wFndQLqU1ODCsjkElW24OduECp2LPsnk34kQ+GLN41oDtlmR/Fp8UdRmKuIMC
u4qDYH3xwpGm93XMnYUUuFUEAqFm9Q3Ffjhz8MYIypKTPpUz6cmJh5ASPsyk4A774mQitVUNb4BO
oHNa6iLvtVu94vIRzdgN1HCroMhmchd20iHT0Ul6H1q5NcCcC1TOGszliZMnEqflT1Kv1QF5uEWe
44MQzHnwwV0VVqzuR7Dm3LILkgfT4looz6+iYKdEIBydNsI859eGpkO1SnxDSIUBtpgBThKgUEl1
+P6vSQ2HEDqEiPLVm+ZM2+IKfn0Z0/XM9Rl0CQLaPQJlAUwr77YbytC3AImSFpVvHLoUsejndnRF
0/hgFMWSO0Fj88hPBHRl54ctihHbzMIP6VZfd/CHhIKM4kPZBU7icSpzjRbM4cD905RM22OEkKat
gvwxLmdVG6Pzwaa2Y2T+IxiaQ2Du5QistGtBUZMZjWCVMtuaRNoiVBfzJujI+DZ/9D+I12g3puAZ
5Mz7yeK3kSRT4dUn74wR4ktbwH7oTOcVCqKlk+I6jiiqGxwHTzSPJOn/x4RpRJZcLNZIEQvZpCbT
94+6y6PlYYywY+0SRcBVarRb2xKD/xta7QyfxnyBeEm821uM22X3XdhNfS0JppcdhpbJm6UVnq1G
eRoVoNWqRSaixvWgH3tH110pvWIToL6pCTRbXIAf27L1OQSNqv2YlccaNDo8wjnz8vOEon9Uff62
3ovbRBNdFhdc/xbUaCyxtjNhhaKWDiL2BS4cWvmyyDkZtSqbE9PjN7uO3KcYTSZLty0g8xfupkzb
SEzJho3DPjgsWVmjltH3WTl9fcPGFozfLTDE4dNVM2FA7hTQzPlH+4+AghzTIecf2fCTfTMP24uV
jbmh7orIG8qcB50pNtQlyXpgZDfvC2G/w5D/CUmtsPvpOD0u6UYnLBbz8duag+xzTMx8LB4SXM64
gZOhFw1MIcT9goXpROdYvCPtVT16BgmgzN9SaF7KHlYxeS1dMp32+o40TWZRQnOogsw/nx/2cR2/
ksixU/q91+6PP/PQzYFM/BSZmvxeE5fZFZxtQyJ9MYSJ1Zi+TBA6QEGW7OuZBLtPg8PG4zRQr9G0
6wv2Hpy9gYaPef9L5/qi2cUtI7V5c4uQGvqh9WMVys0AfgEyz0d2DFxvyclvD93Stgu/EsgY22af
cDtcxGW2uuytuyKXjv59/Ogde35iFj7e/fLm6B1wZ8TEKAaRM5N/LPN0GdC8TjBNg1dg8uVndIZf
1gHEodRkUh/QT6K6pYt9dExUt5iyK/AREC4z5rolcfHDwfJx7izuNeaYKiRLipQwuGTG9/ZGh4HK
PXsuKIBrzcDelN1QZiMIc6CHmDM9qySFxCowlGmrqTqDc74yMGqQUqQAhLMjRiWe5zoFIvFhgocN
FEClbk5cw+LNYjgAcKLHQ0YpLGn4vCKqSsUQtQ5zWdBcYCyCwE02R9gpK8AL7YVeOBMxbsjDvge1
DOG+waKp/DS6hbJKuzPSfIGYu7ct+YLEOPY8wGICWpeVUAjRITvk0c7dIuiChB+qQYIS5Fb75Yhw
P6PuF1/3XP9FjRZS3OdVddwALivI0Amoj6uj4FB2dF/qe6CH0XYR0cNv21EBBj/9LeO3OYwhqgxm
NHWzuKi1EeN6qc3BLB0VFWfMHNSbUdNVI9u4gjvUSGa6aT2Xg6eNJG/7+w+U8cZcy4v6bpjEk14b
W9ylt5sGkbtVdfM8zQAz4mVcp/iOyJOOH26DK5CIfFkDifX+iIugcmBf+1gVGjrIh3d3k8FuqVdU
IHi490EcV33U2/vc8+98Dg9znX/YKQlPj3PeUuFfm+vc5NWSAiGKheOjDD0YlBwaAbvnt0EPQpcp
BECZ7KM2dSJ/eufDsKSOTdz0o4TqTLB3SXNDdxL33Glmb1PWtO+eH4cgOFm5DTkmeuErYy6ctj1y
XUF9hBg/UvGnLbiRm/rkMe5T/wIAPS6zvaAYNF1bv2U6nYdzElsoFuonx+vuyMiuCUfPxi2GHU1F
P22mA4ToVCUhazOrWKe/toMojKmJTcPjBlx7Q5KOvNuAyJ49Y+w+3tyn8bQFXHekg4YEJ1ptgqPr
Y6motjaK/RB90W4xg1C8tXDqxj9mYmHXo4VLptOlgsNWWoyq12JZWkY2bcvKwYi3MPr2U8hAJlwI
hCGSe2egGCa/Q5mWq768khGzMkb8VrS6ULT0ubo/YOSpecEth8TXSbUylm8pFr/kPkX5GSeJqOa3
7foEdvcwdTDbTnifaWbvagzg4OX5q0KUQ/47Y3tGQ5qxuaNudcXWNf9Mq+fhD1joo6fZAK1jB9cS
xG22YN6fFLjqHZiZvW0H+DepsdA2UIFi04ize3wwwMTGtnxNFEJSX02kuqe32X3nA5eVXmygzZmQ
2b3MBJEW3dxeKvbmAC9UpET4eirOR9gzzKb2zHB41U+A946/8GHxi4tQR8Y/2BnIARV3qY2hNl7K
XzcFCaDDa4mJZGglOvUeSZ0gKQD9zc4IL2maiOg4s2QviI2HHkgNwpmK3A38T/8mBDzQ2AvbYeNi
K1Dv2rf/jqyHdX5TLVabiYM7DKCCfdiJwcRu8a9m0NTNKq7cDm8VLXatayzeV2sAuqck/veB9uQx
4iuA6yIdIJz+oQlIgUa3P78WbTb8ExQ0picCipD+bhjoGI7wT7S7hRxF1wcwfWo11LpDCPVxe5PA
kKW5D5/qEe03okg79xDTMJ1EGe+nfqxYr/34mbFumen6iF4SjlPY77QsluV+e3dlcEp+RkJ8zw+I
Fr9jDrvyQa5kL8DfowLbJinTJa5WOAAzdQFJoWM8IKA8mMuPIIKBvuiA/sR9TbZSegNGntlx19Nw
fZKFCS4KhiGtnt7VWdCgRoeJH+XvzDQ56+IXVJuldEnYey5rCnnUKIg0odi1lRbR8CszFC68q6+S
DssWvbLhHYv3JwkgkR5vk3OWqll9Z5PtHNR36qQLckcHka3pbF8PZOc2cfy8RqupUw216l6M6Ynr
+Ozrjyr7iJPTeF4ABtCWVNWNyD5zxmo3MOIRxEUnPwC2FCqurcnR4L1nsvEIkIRhWRWPiwFB8z7r
i4B9hHGms1GtbZ/D+yFB8oYkklPx8K6w2YNEv0d3YCPpyOv+L3oTyN3fMnf1dxEQ2/kxlPEGaW6H
P9+yyct5azDaCGLjs9ep3PB5UbDYyE07iS3Ji8HrxxPqdyDV9itOZMv6oJvN6yENyB+UhChWE5DC
mtxNeJj/O8tWZpciaJC9b85V673xFU1SHhE3RXh87rdKmIktnxzfcD6Zalg+xAdict1w+wRm5X6v
1hQJKaLwUZYecghxYyMXtyaAaL6bIwz6UQzDVlYSTKsbtO5AWLLWwY4FPUboRqUwWYR4GyF56TOP
PpSIKy5Wr0qGcXwA1bOCD18/dgVLy2xDDDNffxzU+9EuUimTQxsnQY3OJkmRbcolIKeVevotziEd
lGO2hseP6sJ8TU/CnTNftnTADNWqMmuBiZDBn7wN1tImrwJMsL+i/HNWQvyMTRUR/zeXNgQ/WZlq
ZyGR931UYHmJpmw0rGKEsXEFvndVd7oeRgi5YTVOVxmaWYpr+C3zQ7oH93MTg/uqoU2BVIoDUrcC
mDdmVYfvzTeDgxbkK8CWIo9FC4rrZoFlcoF9cVC7RdnvJ6LXP7G2OoRNQL2FdQrQp3kBwKLaY0VK
1WCxKtagWr9WVHm500CQnFni4/hhg3dIB1uL5pNMod/+1FRZfqOcVlHNoupSbYn9TjD/3Mjf771r
bMDWVE0K3gQuNOsgCWiCmQKM2M4fikbR+yJxcN2TWYMIftUcQneA6BSymUbpJKIgLBO0uDoNEV2p
KejwyfVCvN6jA5Et08KQTopdD/5EfpHCq/BVuVMOvVAetsTRRvrpLSqmuE5TEJcAeDNryx+TOnyv
RRC/U7Ycwz2TJSm0y9/etLOWMyNaVJrv4kbc9IxNSEN14S33P7GjvOHsekgHTRU5rCiQ1o+aP8hF
04+T2pooH1Z4u7WlRjktKgNY0j9yfvXYfOGqJ893ruizh0BIeAtd4eoF2rvlAiGMgLZrQ2UlG7+u
gsuXEeDic1vuGT0jU8CGUNzzoWgryAuvEtcNnmQtztS1e5HhbNxqpekYYfNG3iM5I3ihkBYpa/cZ
PKQxg+7rnJhD4zjPLLZ0O+0lx+CDPXIWoH0NAKXxnmYbctoYUA5NbN9ef2qVZ57sE6gx3ANBeYCT
fMidzw0MXE6XbG6t8kB4IBFY5r5pSsO8aqFj1ia/blbdVlMeAzooS4nwhojT12e6opg4NmnoLdOb
Thozdn8LepkgzqtHiW87qwCjvTph5PklH2QWBbs9FQ7IO5hcCsm5W3sU5pqOxWgzemjJ9NfkkR0v
PWsRUZkp1ImmLqCByJL5rzHc+Qf5O8zqqeSEiADQoWJbCF12bC1DxojRIU+suSMdTHdtqt881uKv
9lwbgkqXlLfoqrpD2cZ4nX/ZizEP17ed/iGCuBODllDu82+F3tGrFPqKFEu+hgmXPYYZ463GN6Hl
IawiUgLWKKKB9pm8U8xAu64G8uR9cX2nRCm3p+ROyqv9TF1YJkNAbSneGJkf4SRG/pNh2xmVL8Ij
5V1ygnpav2PFL7QdH9e7AHXMjBn0OlX8ZjA/+cVcqDBBiwceAXcXsbAsnFXCKzGrAdz/PiBUNPIE
h4iPqfuyfH3UK1lWZVWFOi/QhU7mHiWDeS1fQJENGMyYkBuiJli90qWuWXkw8d75hK+zo//tQCcr
oT6DlLMqKy8IM7gU7QXG9BlAnVlXAiqqM9lAgUpkORabgF8a8AY5dnQwkxhexoh+0ZJ+NKT8D5O0
wVh66dK7AJ32wKN6hiBWxlT1z6G4219eSN2+2hsgnvDBhkuShw27z4MeQ3YY+baFlVrdnTu9TC6P
0AL0zoRRrbKlaCPBgLh2W3RJn6ueLzhW4+FYPD8OJbUkYteGezFRPw3XE7rTpBVP+ENy8WsrPkCW
wlAgr3XV+pY0A4no7idT0fGPkE2m77kmrzgUNaCAuhwdO3xr0s/v1zVA5evxtNSGEl7N+6bxREJE
7kOt02PzdgzgoLbTrgw3n3tmkeiTMZg+JtVmjYTO7XvsZaaVP6fMoogrsU81TLCeTfYbvhQkVqSO
yFkrnOtmlRskEqFIGcgjgw/xkb3O5b47IBE3vx4kEOnkX7eDZ6DXhLObuLgkHmIjo06wi5oJpArh
kqLtZY41p+BiLgm8OgOVTRvAvY8x0l9pkJNDtJ16M3/lE5uLiuYGxX+n0f2UymV98OKHSPgixOPf
deQktZ5PxZMP8AGk1nUHv0geEwtFyhBhxtu7shFFKiQWJxFxTEvmJIC0zCvRFX5tUp8vxSITII5J
NZLA5x3yMSb7a9GiN28tpvs98ENfEJ4kjrRxML9F1dRDxLYQzMFjO6DCmsnKOqcviFQ5uYCbotyl
CMNooIu9f7t9mW9smwsymmIpMesffmEbjYF+OdF4olxe2qpWjIQy5uT1s9ejz1F69T8/gjogF7uZ
kCNBwrxxyqwoymV3tFrF151f3GbHZCvE1DZuHMllYJkE9oWTeBaR4RWjj0lo+BTyaXJ/7iShrc0C
wrV6DlT8SnfpcsBFzqYuB/6VV+kF+yoOILVgxGdA7RaccCoH4BiZ4scqGdTyenUwSbdXJyclbZqD
DzwpgGIx+uCuPVzLYphpbgeDyJPnNoP4uJa41WZdwssxwtoDx+ru18vRAwLWF54nvkj3sKEGTOiv
9VnD56SUUoqFnTo+RjicaisKSwf5Omyuns05TyAokTB+mV0uieh0zlH1U33yeWjZ5RkWQlxvx9et
R0vtnyMU+3T7OIOEdpjdSI1NkXrFE1RklaURqzsKWM04Z2s+JVJ2QZXb0uj4zxn1p+6I6OdKTFmh
+UcdjnnXx9GtdsK5uFr43R+go1t1SeSbfqa0bYTT63M6hMOEthHXOFxqfk5stiI5RUUsmN9PAtXD
e3Nyje2BncWI1MoAScE2E4/irXtqz+SDjXDKd5ZoKKLFZc/1S0jwH4KHJs8Ic4fLIaz8462yq3oF
rt++UIImxQnxxlYBOrpUTRJyV/uD36Nc2pGrh9haDTWmRarqJfgoFn8dBqCIe0oOB8fLn3L95q42
wVy3+uMHW+d326lYQUqjgKYTZbvw4nylVh7pZgv+D3zMVKXceP2JekaIUn4QYLxe+32zZA+u5zNl
fS4P935Ww4LXxdJH/M5qlbWbhrGwazW11wsfsS58OO5r8zani3vI9NnnP/zwNsJoyyaEHn8JM0/z
IbiIpRaxpsgPr71hsKKq/PRB59ZqtTkNAzlLiYyiWmcgYopGAFyZQ0FpNN0+szG8EL4IbdcnaKDb
3vUw0Mf6grnvVnYo7vaj+ZNm7aN1xp1sueH0gyv92gOFH6wLEDxNdLNWCASO8qXW5UUF6s7uDpvR
hHyaay6CxpJ1ntdIdYUv7RCe6X++2d62YM90h2+eu5hrmn7M/aIVyS8R3+Q2zt1K5l0A/8NjUkzw
EuM/Y/ZwlRkhyiVhlpXde6zk1KOE4PIePxlB2USN1BOkhTZrlKS7Kk9HPQzdWJvHi2GCTVotWVQ4
Mx3g/Bjzq48TZNKnXRK9Uy+l4VvYncvqqtHDYJltlRcCUBvhycPDBPNebLYJyXu23TFSiBszhlqc
XKMLUEV/+vndEc9u2d/tYLk8HkfW8nWIUIkCegcHIVXLh+s5iWrdsDH1mIMefzHQDbhjz94gfxec
2QB1nY5GmqfzOS02Zb6HmxXUWulBPgEU66eko+7NnIPM2DwuuT23xm0+7t/CkuFdxv2Tjua4t4z9
3dGb8zfpVxpxmcynAMn2MNS4mPnCGnK8456vuqJkY1Ul2ybhVbGZyZpWrAFBXGEiILDGKYBSHmJ9
4yGL4x9o+y/mGDUqTSo0AWEM2Xt2L4hkVs7gSAIhlt9I2LUGAxx1p5xA49BzLCC0QLDpEULqMebo
zsJCu8KWM5S/zjMSmy9M0H5093baupIJkzcnSxReYGNV1hraofOfUwI6mVE/cs+s1zCa07rT1ids
uFjsd3LwsCxyO8OxdhpKE+JDzNm2O/ruGVJWTD3PedIcSKgexWGogqU162KgR86xCRA4AIQrD8Ug
VxmgI2HDnFtqMBzTxvw2Ajop/AAss0RXASn58egDhlRLRFWOY9vOmSPIDbGUSHEKwhTTcI6QxpMo
6hMnhLc2ZSpjYptUsG9BIF5OnLb9CuY5Ks3TjQE5ixvU8kzrFUDkRHGHfYwfKsfqmRhSJ+rsAyrb
3eyYy8SEmOGxPBWCk5o2k1/Jwj63QOW1BIJ/EwSbuhPiyL0kweFXb1PkEP+A3rrMbpRReDzq4spN
wd4+x42T2+1sCOHLUpnNzDrXYDQHXRzwuYvxO7HYhKcjiVtrpYOawPc+BpG6dLkQ5wL5KBdW+qtD
DHwhi+fIBjktBdf9HFb1Q3ZBAAIagy/MLVn/EFtjmyLv9Wq6FoDTyD0bDoKxVTXphX/dsIaVmGcV
fD1Sl9BUNzIU4azw2K7DMobp75+0YmXZuMthUpiea9b2fN+6vbH5WuGtCIf+KOg0rOdI7sRpFgJq
ZuE14z6TlVk20MaOBsWqzvuu7TTGKj7OrSIkUKXWfPQ6F8pvAQPBCqnZrKq76xQxxMV6Mz8uJ6HX
N4yFkWCp1ojIsGu4y71YqdqM28w3gI+chfk+EeMgJixTOCl6USL/vzP5MQDw4oflnjm5J5zdFugH
YTThgUpFLMC741V/xsliSq6LxHJxdZxamKL1NSoYbhgF34fqtDwSbUCWKJ5JIbXZjb0oOPUKdLYx
VUoA/ojZXhwO9krkUab2acEKH5VjJCY5doEamh5ziP5zwxKMlNHTBZPVkGu38RGZrcj6VZfZx6j3
P5LMSpnTXdTt2h6OlfyQQBWuf403ugsOXmshCaocE2c3LuG5iJFd2ptcVZq4Rie5wkyiEjhJ5nek
HxQ+vrV1pxfeMngsjIOtUOMNoS9HjjlTBegweMWI6J3uNTzn7WgIgGtifHN59ck+KnTCvxNEpciB
4Nwi9dkKztBoMP3o687ErPFiNYkHFsliOMrZzJ1Th7ekyvVnjv0TGzjvgwR7ws7PWlZGN6osZpno
ugKjzDEOsFNJAiJydCFdv6n6+pm07JFTkXP8mxxbZ0z2MsoVh8UW0o3upb9cVU0DhJDBaSTeyjSG
1lmljW9p29zswgTyZ4x9J6L2zAsUn+QTDlkHYdqflYxxyNaKMLGE5uabQS/tlza1guVJxFvItJei
C38BCKDliiLkdXyWuXpo2HmzOmHo1hP1DMB7e1ixGwtqCII1v//sJjgN/NFEft0Q4C8m2xiMXEIs
PaufKWM71ZiihVAHFzdifxX2rfteZvMAeYdJh/BqOCjVSSC53l4KMLykhN37JLb/XpdQX96dn2mH
xor1F6Cqk+50vU2FeforQd5FWYuTpvqoTXOKGdm5T6wMmLI/Yy+63ngi4uPml6rFWaLJyjuWaljS
OeAlo6UpBxnfh559gyIaRY1XceM13OwAeupbQLNT2Xufran7++F7USfpcoKKBHEPxmPFhf+KKbmi
LUfxuhUcsZAN/LO5a0bXuUV+/imrTg/okE5aJgvS+zVas24L7lDw6/eXA0vzMCB3YAceq0NSR+Ug
8IeELtFLxW7Q0NbhX23s/JJysc6gt2XhD94tIIZKNVxrIgnf2GMzUHJPAv9sdAhjl+PcKsRfyarY
ULA2aAJY26XQpCXQM4Ko0Y2M9rnzCBfkohsl7BhhdCYelK2HW1so1jEh2RE25Xm0n5d2r7eAkck8
+Ta7636ZEvctChG6I7mfnyqiqNjKCDbLZOtOUAmv/9YocnFsqvoFJ1gMtnH9N217aBAEVFx4OchV
jMzOuSQJt0g+cNDzuWw1uINRAlej37utI4WWiVMdGibXPXGjuj0hgMK+1ilrKVzjT9BkajF/UjmI
o2DeE72/2H//vze9sFcnULggwazX0dgmDmIZoOvUi3YjVWr7uXBu1iQ6Su+Qo4AyYsUd7OhPpt4E
owbQqEydC9NeZwIE4J7+/L+l3K2gActfgeScXf5DZ6+X5k6hZFmY9z8F06HKiDFXuO517+gu9IA0
3tceKSKL4CNsAQ8akVrwJeP/xgDz/53ngKFvSj4V1Saqk9lrKZ13OkSoauEco+OuTgF/Pr8WgvZ7
CGFBSpuC3hRaZcpLY2v2dtVdedQl+OtwVAJnj7PyW0dCWAWFtEUISuv8jkpui/LUqbWvI/yR8Lab
0D1aKWdZRvzl8VHocDh45YeLQHeFJb4pgGTXtdYwBNKtA/X/r/4b3TrE5ivs2OqNEDKylY2YrwWX
xTXdN/EmVFFOZNFIlHQObur4pIg203eFti8emS0Cii7As+SrnBXVZP2LMshcX336k6piA10fvXdJ
WUCag7D8rADV3UHe0jP9fiw9v6IaCtGqfJRrCPRiLsXrxBaQtaI0egpINksICl9NdKotAay5jrjw
tO9zIetlUrxFn2MjjUyQOQWYPkzk7AJN3DbhmhXS33R4hmDdlwl4w2AokoXUFvKdRYOJTAO8zJ3n
yOnl1D1I423TFnphKcgll98zbNEzg3i2wbN9NzfLOaITjV7BONBaFf5WGAPPHnNEsJPzaPaSKPPx
WGwloxVdFHLPn0N+YGQlWuPV+hH+K+h3St59croRcKfrln2AjtkU/AjolFyDQ2xpaCzUa1Teo/rp
opBe31dVgFKxVJXsPyl17tCXX6TShYuGVcvlk1puujzhWDbmwOOuohS42QMIFZW7PgLsbAbqwzd5
C48tW86RpjF+Ida0Et1DmuvUzN2seYBRsOiSOmis4q9QRFt7jRf/Xgobm1sqEWHjmsuMEXgLhJOU
lXU80vvKyzIRjL+9YAskdKvPK7WMZE6aWnZIp2X91PLkr4X3oatWbjULewTgr6lJ9y0uOL2VRRoC
jc+sIwGKhp7mRKTBk3PZIV/yUxkjOyiHh6f30MJ8l2T3yr2Fxt0tR8BWpIeHE5mX+OvxvcwLHH7Y
FcOZzZur4rAVnJXgAD1Mg3ok3i0R+xDR9siqaPiBEJ+hhWTVk7iPM0jqqlWU8de6mmz6wvFVEhVN
XOkcQlN2DCaEUS24F7HJlFoY93+h68RTCg31uIfaXv5liSZZyGZMMvxaLSjzYEWjkdps58EVwXIU
nQtO+o7jZrVB08cWg0lMzSKlTyboWi+pzs/CGWgmo/ifM4FECdFSGLveYJTTe0JAhXwPiAzWarqU
KOMUfJbXnfzDJvQlvaLDf8tv7Phe0rikH1YPJLaNTLe8HG3cgEVw8bo478D2yuYu2buqHATkIinc
foBw/s4DH10FKth0NsgU6L0QWaIhQ9gtCaxgJTgin9I3FBmBb0w4oQY1GrDow6XKhDP4CRsfhjCg
IgP8rIpwnhcvDZmpiHyDK0acQjmyblNRZMG3LAmCHi1WeI3bNoNZep0wyS2HzkYOFPfLF13yOEjh
Y2vXQf3xbzOEKCSdUVyrjFTlyTT9P63rX1BN5Lp2NzOTta2I+dJ6WLemcl94Cfs47JhONdnRsXWQ
ceYdVRi1smFPyB056cT69wAjHV1M41K/rfRl9cRwpRAOhoouBZ6W9zZ4TvFjFj5nNBakBxWKF8vV
9P6Nhzc0d1AmpITsy7shIH2DsLZfCVfdTEPwKVmA1QD0VPMYCo2KAJEpvhZt4MGzeV7H6zWZ7u+e
+4ZciMTpumXuMwRxQuuYWBO3GnB8R+2SmvnJgi1HnXPSQXDdBB1/eeoewLIZrVLk1s482gjprDBt
F1lQh9uyMqGN7HkyGP5oB/X2tAbnhkU7D/g9ZY2ECHbmSw1Do1amt9Vc9HFEcYtXE2PrT7fC1L2V
pXNa5TNZkDFlhQt5SrS9rRCfg7bQxDyIh8My/8MLFBArZwNVFE5xqN9ZuMyRqxz6SerLBIhKnBIV
Cy2LSal+WW5WD1jdDGyE1vVTwwJ5KD0d2b6wVyx7awlhym+4zYmFR4jfZA0qHMn2Yvg3pl/FMvpl
cDhm1Xmtx1uVQWAfTVp+JjoKa14KiY6mdV5gvyaDofdVKR10YL+Kz02xykJoeVKAPa9yiYTOSKyI
wyvcnIV7TgEApg6u0KPKRSL6nwXGvODIUjjKQ3K6gB7+y7YocS4KYZ3lCbnJ7cyoyX+9wpHhAEe6
zPfuCY1uth9EQ6/9u4EX5at8IuRMSs1n7yvdn+BklJvZm3gY1XadOpGrbav/5rz37/kC7cZG5WD/
+2jWdsYYEX3Q0NwyNI7vUvQvy4NwbAjiAnmz6YZAR3O9R2qqFzfOJt84J16dFGtOQ2yNx8G0FKxo
9uKhoLZeSmbG1Wnb5YWhcA8/jS+ThXYoDZ1d7qfdrUdzD9HWD4kMeo+rGP++ngC6dop03Rg5bGg+
EbFZYynN89pIjJn6LyS0zG51XdLypYeUXVba/hDypdOJFyBkUY2bTIzJgdMXub8XmsS9zECJuYTx
wti69VPwfZ3QBBDZ85dLIXps/3s3mRY1g0TlRWhi8xt1D50ibF33Rx2C09ePmG4XppzkSvdRZIQ9
LcdtXFgkvFvYJf+QL0XbI4Q2frkQldtZUsICw73cCCeMCnjERR8xzcAd6uvwP43mquJpJEE+Cfqc
54cQutjy4VdUum47Esk3teNHOWYNdbg7x9swQ1gnqdqVeDd8YlIhdATAIp5zkjQvke5pWHqWVHBT
MdOAj4k4mlzwPwMvQ8MO8pw+Sy975NMV2iP4qEmjBi2OPibrF4lFEikttCbgcykJyl8G0OoWtUpQ
py2IWQ6k/esIQNMnvgiW1cGLIkqm3jopaZaohRBptoemVRQy/9vBDE0oaxKCTzJYSx/6dVE2IYig
5XyHvm5wg/gc6OuqOEaZUqMgMg/BQF0iItPCqu0y0tmxenP0Pf22bnXEOS78EFoUdC9UxFlHLbKo
pPo1i/fgblC7uEgN82IQi5+w6AJMJoiwJdkhE0SbYjZAdBaII3gZuf2pP3X2R3ClnkqLwX0Pspdd
Vzr+uOvnPZLqDxi2p4SzTbLJNuqPvQdC99+KPdLe9Y1P1UdCrQQX0/rq+/mgEcAvnbu+vAdIL7io
sUJAIX2jOyabKMCzreadsV6XCjXGQkk4ejiKljHFgYPiUV0E1LmkcHvvW2dc90jcN4c8ykVfDz+X
58YCXFRaaCialu7YlYSiLQlSLE2ahkvkgPPJlTeULPJjgLdE0fk1WHcPR4i37HxDfEKWlg1n57UC
IgSNROYAyo8mo3N7Sl8DNTAnG83SjarwO5h+TkLNqLdV/Bj5odmQb9owVP5KoezWuO/VIq47ONbB
xYoBzxhyYr1jGo5m435hrTdM75BsEbpfHrUuz3WNAlzbs3NZ4zhH8YWoz2OFhW8Ov1E/DPUu5qEq
JMcYZOT1yYYmiLU19jwZeS2gOd15xElu+V1uPTgLtva4BCgESDHASCS2mHOq24SPUJNzX9PDp7O1
AOobclOt6b1PSeAO3KwpBjSBMdrpdjF3ZuLf4xE/+I3ghyaCc5NcfUfYMEi7/20Y3JDkh118sseR
5rkdLMPWUNhHGUBPdh7aciAX5IT77hs/xFYHp7m3pUVjgEH68+iL6MsRMkyUCf9c9cAHTnDw0BYr
ewxHXZMbTSsPy5KLFwjiB5PMBnUpM2O6j2NMqPz7XgudWWwoi1rGBXQkqE1OBGXp+wkAsERWtmxL
pwyx7LRVEhG7tVfZKA+07TgDAdFj6DbGP9bHdemD3t3wNERZEgW2ZnE5YtEZlWYhKA1xFx0EKlyv
VhXR9GMXoZQFJRA2XPWMmzXwdJNfOlXWaoXJJY141ohFuPfGKk1d2QdqmgEfza2lDTzcQiinYuio
2DwZTF8SCz4IXoYvAha+p1ivQJmQGH2DtVw1S9n/0MsiRv6mnhGRkuaefPvXd+v+jxE/lYLFdC6o
I9zIgKW9WZ0FzZTxacixbZ7BNLz4E4j1Y+ZPHxHApK12nCxYF+UxTyrXTphOCyJ0Piz21Bof730v
weqKlWy9LUfT5jkYm04HLiyTCN/I1uPQERSk+aKyjSYA6NpU8tijzIagW5LOaUInJGjXUa2cY+Pk
0VCx6F7RlCXDVQKdlEcS5Wp4IzUQMo4MdhTJh1kmyg8v9sEQrmK9wzm9pduP6FHbFoLaGy03mmKT
+oyEWFoQnXrCwHfuW38P1Mm0cI4cDdWKnO3Zz8i8bsh2giNhgjyBolGvNhTg2JmaSgpn443L6QOW
xW/mY4XHNWUQZF4oRU1xLxQf6lJRkVXbWG1CLx0HJXYvqXNzXgHZpuXbwDgVznD9lhLdeL6Gh3eX
AUGXfAdmKNV4rjHtFP8b832QaOcnLU2zJYMAZwX0pZKp4M0xzzJQqxhzuHkdVQGA83Vhydir1cLq
8ONYC4dKH4sZIXTWukz/9odsyXLl1ZAmY/fE1mfrqpyTB91orJZyj6k05mZk1LNHgPo8mIdfJv1z
thKObN61lLBczQM1MTA2kHqO5DPiHaEnjnYBVRtYls2szraQJW1etdx8zXqsoJi7fXRm73YESFSu
IDE6ZKV87xzSk3kTxngf5GaOUrahJXtz8RSObLEB7hlcZAckoeg2uAy9EdNDXYp88CaxcmO1dTTx
Kh21v/MlX3BOOp3OQNs85jdn4GV1fA8sYubHzBOyUvXfSsBSwODs7TftB0UQUmrBDo6JfO1U0IDY
qudbicW/CEPRKn/d/AiCiHZez0C8pXOZjy43C06el8QJ2o+D+m/GsxG5kfuQ9lpUsHvyezSQcbTH
7dzyPHfvYJKyJJ5aYd5lH50hGuGVIqnIvnsGR+VaqT3yTmBl7Vokc7ZcIY8nPA2R2wNnP9nP8MPz
nkBstFAsJvyPTfn4nhQdRvOmUrFC4ktkd6T3/AZWkwIrWWZloL3oaMfifKueqA78pdNj3DTeCMjV
0eQm7yCh4hjmiYVYTeIo9RHXMG2zbIeKdPgaGC3DrLSuQlyTKiiWafc6aGGhse0pWEMeHMJwC4kY
fQDoDeiyvqtO506c0KOzotX75qdao89lPqiVn+DAM+JZBZLvtdVyZcKPwYx6Ycu3nJVXWZ0DZBPi
yisbS24v8UvkSSQOobq+hkiH9RAxNMWUPGdbOfLbkcEhDwP+9D0bP0a8WTwjXyG/tt9MED8wkwDU
ANqwMfum6pAsZKV4EpjBRi3fbPl8VL3qxaxAVuV7+nyjj9g6OqIf4ELvngYGjOM8B+aoj8RTXGqR
8H7jbzfgKd+wQmDTEHHOLhO4+DuLTLfyTq4PSntM0Vv6fj87pf3kKiqsMqk79tz1wZUuZU3IdoVH
Q3TEdmN0mHUnZ2ZXpmPKCSQv6y7sJ7BuWuJOAApXjSPVfdWTBh5Qz7IP/t7lpnZCubAYuELffPwf
7Al4o8HmT3dutxIb02nvShJofWcXGltKFeVWM3q/C1QY0XvGIkQ79DXWK7gUb7NMA2USo28+1s+7
fZVe8lKm8U2dVwsW3dkqIeFbJOkmtKbPAglszE4TvvDsGxJVw3Gvcg86wO3dMjqG1UoED+AWGhVF
v3GrxaCkzRpS5YYkerGA5ZxnQum4xeofwlzl0bD5ySYN35ScJEgnvRgTKAXtcgRquD5Rs+AXPNrL
J8AdGKLftdU/CbzXM6hGuI3dsr8eHVBlOYqn7dm4+70+h/b7HuKpybuILtFLjXO9mU0zLU8P9mVK
nInyUZrqZyj+mSs7PC385pM5SC6R5q+jPfSUVc6BEt4oKlz1mDcqrC4hnGAXTB+9Mq7A+0/pV+PA
vMMpGw13Ec4o+uP09/Snwbyk5Qgk1xxsPQa55M2y41xhCAPqe8W/uq4IU5IYSzuIH0kNQkDMPxFS
t2xPaEPnY6gR6HnT2jCe+Pv6dFworRGUXB0R29JUt5+BdLjaDsTkJuOobueoTMGCdhe3S2p8xhHx
BwMmh7oThemt5XoVnp/sHp4RFR1knNed2hmF14gx/45xD8cL2DaJaHTfY73esHeorPqvSIfY9Td+
bfYbBas/D5ckrzvW+H2rHE+jPr1qYkvnAawpjLlBPiJQdQlc/0tpSsuKw3K79LCm+403enrINBAW
qztnCH6c/bydzxHt/NeMtNh2YBuk2DUlPyRkZlNPmKASM1UqqFvjy0/32gR/z36kGCVUwAju9Uex
pqx53x9qR2dyHmOtUL7LPq9srjkPclDq6USJersIpbboodNYk9AfC54lW41L5F2ZmREBqI0yu7UZ
WgkeJfMk/a4LBMft+8XwUnoN9dJffAdcHZgMZdhZC9oK9O9FGFRTEkprxDJ94hzYl1V7fnTvS+3l
bvCvSrBtpAfYBIn0YDyPKD2gSK3zY66L8X+Ia+BoDM3wBgG1HYbtxUhRGS18TpttqIWHyt/IlLGP
5ky++9476rlaX+vXn0epQNfK3yULoGCIkJpG2O7Owr+KnoePL08Ck8w6cnSbR6mJbqhpgemSNnr7
pWj7Ymty2RjI0GSKZ3a2kwsPzWLNfajWX664AEk0pYmbGLXR+akXUUSxJGQLpJGOSANbz7B/VxaR
aevZ879azKC/2TPiPO/8a837Nl799fRWrK8sk+2FpA6JFXOw+zOj1FAJnDy7yET/DtPS8migwDXY
khIDaz5aPE2icJHtOpsxacWcEsNm4s65uH4NGTIiA4f8PRvskynmDO9Pj4h+1sWHCDW+/rgcFaU+
dbncCTX8mG7/pYpwNsxVxYTEZxwwxD9dKWHdWR1Con7CSGcMxAZ6JNGxalg5DJt50SbpDELj5zuA
KAyqYdguVUESg9iDdTtPFrsSzTDgDYqxRKywcvex8viX96ncihTUH6GwENiwoSnvdsWxN+l6NcjA
Bf2boqMj/UdlqzGWJOhmy2zLTQGcXuYqzBCWVsLroVU6+SYQdP6Hf0mjUHkZEA5gipAC250te6QW
QHBYMIZFZfOCVHgelZJuD0fVig3LXavxvroVx//GvhbY331GTNqUh8c0ZFIpaWy3aRf0eDanzasy
hCCFHd4A4BlqPWyLO+6VlQnapEcZc7iua0sPwmTbTwvuq0p12ANn5HFAlkwRR3fAPBCUJjagg1lW
P46M570RC9/6LVmmWHbj82KamC01M/l0E7IyHG2sA1G3zWsOvKlYqVREVULZ2T3Ala2fDCG3ZTH9
T+mvM/RLG41frgYsUCxNugGEu/5b5f7Bnq+0S4I2Y4K4u7rG0lJm6pK6IGiswwv0DC7htEuYbwF9
qVUwq0UGn5N0AV61q8PNwEHVw6LQtAyOoZKhHziUT6jAFjUh+oF9FmsWw0jV06GgIdAgZ+AHnf/i
WVUPZTQ8X/MoRpnFyt2FpZLCrHhN55FyIE1TEqT2Tfl0x/LWXRc/fw/PoJ5J4f20WN+pf1cXMoNK
ekR44+Kp58VX9AmhkVCXJr5MUkVc11j/32hK7cNzSyrsZvMjAQsMazXWpFQ1Qxu5JotZDskoDwKf
m0geJvZopGkY0Fl6Ccc8jD5UxwJT3iCTHOiS1s4HyDV6ZT/Kt70tiCg4HtW7mhmNFngoWGPN3S16
Qb91duVm+48Gv9Qowa8MYtYYw+wG7YoQEe2ptIXCnyh9/YZxvnptEDpTKGIuYDy5rgX06wo8xZwi
+yIOVLC3mjV4vExzqAVojmaH3sYaDIj8edYXO0JvgIhVAPpS9axgo4N3N2azxT2NzguZLTOQyvco
tIoGTrTtOFfHNdYvsljfTbs/3fGbd6QYoJcZ8w2JttagcHTBdrEKiNx5sNuMS0LjRXyLjJMzX6cq
lImTmmYEtBAiAFUYbXDIWTa9Rz/qqfTpihAiL82MXfFldDu3thCFm08bHndKoQ1iyBupAjeaeI4i
w/m7SGXg8OwZhDklYO/MjLri0RtYaNdIaP9PPzrIzGUzKZtXXHZ2mmaFiqvUJfdTQw1p7xzAWKdk
jHCES8vg6AO0BfSVk8lteCmjkTszGvtYka83qRRlbvsP22OniZ92jiOpT6TpO8VGL4kBtpKzO1Qu
p9MbkDrGZi3TCCd65wFsbNGnMxLqxYgNr+7vuPg/wszi3GcXSQXhx+JrByjiqYghzSYU9W285gr+
qWnlpVLkc4TbTBCKlHtr/T15/mlo+nv07p9v3PDAawKyBnRUi8yBdMxz165qiWOzn0smY5P1mblZ
wwcE3zQQgOoBBYJuj81oK/t8m4mhJeqUsbA5FcMrYL4l8uRqqBHHPd+2+g04Vi4RferWbu5tpRVh
/XMbpzMyMEjGwxKZnNDOQ+z5NSBHY4rHv8liR6HlNwNLifenCxwJ33hxu26efqaCc8FIpC6jnVfK
W9zixFDe11obUKk/fnS4xb6RVUOm9gvUhmL6h5cTAR9efxC7+lIRlR5LlXjwN7VwjfERyB1V+mPl
giNhAztInX0YYdBOL0e23ZfOc9X8X1Hn2k73meWaH2RkbswjNnZXg5TDF2kItQ6jcUSUJEzNdWo6
cE0SDIi4dofyW6UVrqwuhAImx/wbJMIRBX4pVfW06VEZmEw1xsv2fg75S2QoxZadG4+BhF5f8IEc
IE4D2As/G7/6VuCtLYYvrre0TroXu7XkW5XAziikMCB3hj0iiT6KJhS8/ftCdjK3hPoFSUZJWp5A
3lpxFO015ldvIf9KlTegonlL8co3i9B3yLAKFoKf4Ezm3eF8exSHYgUH58pvVXJp8d7ESiMMWFrR
c1vgaoaPahGQvRIxuPitUaHg8I8xKHcjQr4eycnAV8plXPeEzgE46jsUgFYyV2HWV86ybKvrG2Ap
JcDV6E2PvwCV0oZOq3+XMjmXypiiEbfB+/ix9JQlcB/Y5T8pmEL4dOdRWK8pxJRLISkJHhWc83BR
v7B+SxW++EVu/k60kyqDWe8m1JSZL5r6Ycy65ZeXwe0yThtWmGo08fTWq17PUG4hwK1rkCBk0ppj
F2gtdj5AoOjYckwpjadcCwfrVr3z9BL43iWLrB5E4sgKFzIT3ir9XZvOKqsT407dpNHlUolkjK5K
Uk1ysGmQ6vtSN8ovG7c+IGNkAlIm4CHER8e1qJh9qYE2HZzgPzAKmETMlVPkDp9RAm0ALdeZjytT
uT/As+RK7Q1ychdx+NQgI5KwZ+v+Ax51C1TG6BX/5AfDB/80JyRFBsnx46ighU/5BaoW3pAxYbFq
K+WFiQeF0Y0xgXG7DZwSTz7H8hFQUrYauEvUprioyQbg3EyXT7a+vaAuYCfRI1Nm0axepTGKD3Ys
IpkE85P2aF+QMxGkxmN35VS1D/jNtISNZ/ZOP74sqo/sXeM0eP90PmSt5OHxucPrMYM6Z+G6Lidr
f8toVVS8RzTOANPp8VzUehUj8El//+Ll77eEXlpcplmt+kKgx1pR+HZfFZdmDmkiOrMAxvC2xezH
epT5GYKawbXDQGj68PwuKO3wPgKpkiElXNikwZzep3xEEKTKlroXBDoZFToZ5skqPgpkOI4QhCio
ybBJk2B8MDflFqMc8NR0NYUhm68XY0UQcinc1xRQlfpfdEY5sjah1uxxVBAQRC65XooCYHKbf4PT
EbXvZlgG9hQSWE9nitXBXb6MSa9+EbYiTyqRwi0/hWgmC/u1gqUx2WZTEBpGY4EkpaF/1d/8ArXz
ns7oiSbjyfRVEpQT2jU971+rSh95s5aYHbO+AlnGWNdrw+q7v1yFwyvB8kc70BZ/afnMd1MlEQul
82pLeF5v8gm8QlbziQX4hPT+DJLZs0UUMfEP1zE01TJRfW+OuF1vPXe8Hb8KiFnqHrx2SqNWw26c
Thd9r8QSKf3IJz7w5ji7v1VtlYhjveg6ihjDvbbU7IPDD1FkMSz7HJmUcvCj9MeuIzX47/qH12GG
8I9Wh9OwbFt+YaSw2qXLtDK9zqUwv5e0ETLabfLSiFgYmbt6UxMG5foF5q7AbSRT+O+Lvv+jPW7r
35vNClfU6fP0J78naQOP0yCqyosUOVfDKTTRphpa4zIcGeNOggDyHK1hI7FoXJipG7jfU17j9uYF
e24q9c/TNAZCZxgh/ZXYZ+L1r93hTMpM1RUwaypUsu8b5UwVub38xJC4uqFo0xftwidVxCMPgwYK
jJZvVhjLG8x8S199++628MYa5piZCjWH098TPkpSHP5c4CGorAMlZjkH/bboS7j/xkrMLFNs8tpn
6rduomL4lgCxIbuiCHk5JpSFrBxzybEQOEvCg177bnIThqoCcxv1snSobseEz0Ij5KdaTzLihgZT
m/ndY8xirq7JcVJV+oLQKQimZSKJiGqVDaKhenJYiHIfEvwqWKPRUY9fo2XyaZuWepdom2QB6fe9
yn4hj9bHntHuDnXtNEIXnmVChLw6Z15J/eClQ7eiLcIrO7TYml5UUAq9Tm7o9cRBmKP0X6ULWghM
G1DiPsRuLZlPIbRi8dc5Istznzf2ga6wcR4Cqn5hGVBH4zpLuxHeBZehRD0kFcqk2J01XPPBauzR
4fmnkD08lOimzTXgl14Ft00CA3uWWIigeRzLDGjkZ77kROcaJvONotzMVHS1wYguPWtzrQyhpUzL
m15vwPuKpvx7UsA4T2TvqeY1xfb/35kCLVW+/bDaA90fbVM6gPqdwf5CNIAMtnbD3mbBVAIIdDc0
XX7IMAB+l1Bmxq2kYVxpXLZ0/haZNSdu55qi9gbnmMZb9oUL4oP1tueDeCte/O+71gFSV4erPLuC
U+0E/IVhIJKUcLwVwT4qTgTUMsDfOu2Fz1Fe3a7kphip2WKnPJYbMn5DBgG/54pQ5pKsQI5h4z1G
XHassiGLJFXgmvbh/CsRv5uAfl/25MU/DLpGyKp12txyBBZXaZo5lzRYw7cgHjx/vHII2h2r1tY9
6vo25hK3ZKe1Icdebc5jcRj0x3F7oxGDd3Abt9Li9wbynVgAkBtsB7gO4GFb2pc8gZBWLb/v7pek
C12gEzErbflbEX0qyG3Dv+0QQpxYR5pPoGLWZ+rxkaF2tQqwGppprLmvqB5r2b2ASIWSofai0gG+
dOV29KWqCr5lZUkJyiFwhM8U/aGMhVEv4y4brp+j8Aypxq+pdBIzKD9OydhpnQz2HN2+sDIxH0o3
px+4RrUsRc6XSeSNKY2BFNba4l678s2VSTq4eWMHjvWQIJhmcrzuCrwKUaslNYdDQFqdEtjoutP+
uqvarN9Vmw70UnRbZZcgqRhOJj6XuteCtV9dFnVBu6Yqlq72C/Y4Xby8Mnkwoh9/eiliwGbYASjV
Nm8I/D+jQtbBY1mn5eL70YzbRpRiYNKMsAskO9kpNOxkD2HPwR7zXJS4Yg+q3vSDK4XmOGsv8PHB
fyvf5OcF47kBzaurDhPAc/SvR/tyBblRaezDGgWRDIZs2rYstayKjiplHMhpW9+2iFMoHb/V05co
g19b2ZF1DCBY1oU2C2CL04RNlAZO0O53B7iAhrtI/RTOwuM2mIDg6wT+vtreCq8FuwjHRLbqJ2I3
eWtTbaMQy9BBMMAeue+7Ozv6Hg/rmhT4KbsnnQJCPrwrZUf62U09VTr7TPuU9MoHRw3j9kuiOvBJ
2L5UGnxo80Y3So6yyE+qwsYA89nKW5MJQ1lrQlRlBrj5pXqcKEtHHIg4sGvKkunNMXo5lfQb1R0h
AWbzP11P2xGj/83U/4U7itQBdD8mOofzkW318UzWlv88VWqdVgD96EhXll6cGG/wikXhtsP54fpG
pLlDynelblYn9pA7jPjY7BXRPfLSHYmdbSr1LWL5szgAgoodRUv2nXWpDBgyMiyyadiK2jA56445
x34zlvpFwBHrEVzRcXmV0NF09SRC6kPY2T4Qk7+HmOVuxT4TacLxJLN3fF7Epl5tKPf449jZo7dE
J9czPdAhkMPhdJtpTr2f7wpy3KI7evk8qFQ4tla9ozQrewRXRec5SB6b4ewsMSnfZHOMyE3JBd0E
klzSZVpSBoHTPDWxEB66ABufCdmPnslFvDNnxwVaN9lk7DU8qjiHzMDHsRHBke9hr2qve1rovubW
xmfqrTn1/kJ+kyvKcWv1vqPrTtVu0/Syrhv7Te4uAtqnaEf4hxY2MYrprqAh86zMV4l7RgKH1hbv
h7vg++zsG4y3WrDd7N7nNFIwoazZDYTT5617Ui62kZViihHxM4yvHL1ry4f2hbEHTiZKUNZDrEkm
PQCRiDi3/w6vhRom0MokahvabpY0eTsLZE39eZ+Ix94a21FsFXAh3WAOzwBScjhO1xuQvQ5fNzGQ
8al3yLtRgkY+ZhbZivG/KTak9eg9yztusmaYzeBjsSDVZEbpB/YzHmM0okuQg0XmpyhBOUu5+Ea9
yHU+Az/r4dgebmnzbs/DNpVJldTauL/XW1zTqjDyYdz60jZ6UJL1VGmVoPx4BtwlR8SraLqKnctd
P7saZHcJxuxIjusgxjFoqs2dLeNtPS56/Y6cpen0BT1xFe54np8H5C23Bb+kko7+HKq6gNDkzLiT
kBrkDYS/f3Gt8wsLm+qdZuwW2RNxJQjolcbbrg7XtMCN1SNCw4z1U7tSKwH6IU9lsZsB7ljs76/C
g6VOhRK2PnIl4I+PsXq6ErqPBFt54x/xPiW+oVbb82cF47vA06gRjlf6Tp0n1hQSjnGRvrkMdx2Y
pEKO+LdS0wvTFTSQtG8mSDUGnazaWzkNyzAHYcdLlILZc1qdyY4mRUxtTkhMRPPeo4HplkbMiYIA
dvSM1h/5+/MhAWT9SOvnvnYxRSOOqVWTzAgjAFdjbU0oaFUYeExPyVaDl8kNP/rbD1eCBS+YDjsq
rU6JAmLfOfZ0CEtpKkUN5pJGj3bCMESwY+kRZNEKm7FcYhs8qjQ084F6efFAt2oUgSsrWdUHlEo1
tjg1vNB97maIJDNYo7nF3Js1zZ8QIFKFN+R8jppIyHV+ZhJIDV0NjYE9/3RIfbCOjVduL+cM2pK+
TFY7eVoeNqK/O4kQaZu6iveu7tzNCIHewnUDc7Yp1IZgZzw/MAmaopGtjLp7YMgZN/KlU9N/wkdj
xNzlo5SevgX1jsq2J//DIRHz9iDOAW6l8pSarczDS/tSmH7spoUZ57FS10LdaM2j1gaMqkGliFb0
pe3Y9YQ2Lr1gbfmLoyGON9wh42j6flbEPI/uJDCYb1HIwbGesaavr9f5lnvOQj0fZuJnOLi/Xgi+
kraoqyL+fcKTFUCehOtE82syvHtb3etMjTRp0bReAcgB1SQfvgSk/RuCbz5GF5iuO65OVEcxbPjl
T7RuAGzXJ9UG85jKVvA4Mdqk+zBzPujNJzCR84fs4lMtvPOUdnNDIul/W+A6D5vMBML32kt5nBya
oPyCaHxD9tT/6AtlUA7T22jvQmSG/aTIgKNQ5BcsZT6ogAtZ9gW3HFmBpbQdLO77O9Mb7A+Dk0bz
aMQnZZs/md6mhYOQM2k1bykap5xlqVAJdv5ffHIwaGDV6gElCP3fBEqtfolRGwi40XNWDQbpy7JK
KZ8Cf1KzoOUgrXGXPzRD27K6u09dY3WnoD+nsWXmYkVw+H8MPL88uUYfcP3W96g5CFgf2ugdNGxD
A4jiDVEQgFw/YyCS9Uy/hJQyk4q/0cirMA3XMVg5A9AEopcCaKjatzd7bdg7fAxsT2GT4Np/mgnt
ioZOvDYaNXFf/ufjyV23owfzM61Ms0iP+q/cZVG0WROrUYYK5NKF3HfyVgSrkSw6Ck67EsKkTWGP
xWpuyylLLVVXzEEM9wOxeLJlIhvFPOfKTyKUa2jWX7H3ggIfLRWtOcgIfdkVmCMJGWhSOfbcA4W0
eaFG5EEYNrvGRt6hKKamFBez8FO0DVPPe29te0s+vnHIUgDAKYH9QNevSmIkxj7TvbG1sqCYtcXC
pUICk8j5cY7CGDaHiYvA4ZGhhLv62x9r+7No1QPNVkojsbA/QoEV0+Pown21FwOp0PNMFv9nlfSE
tMTR7sm4t11/Q8NQVCeuxHYXfBB4ssTbX3p0qd3xg5kquA+0X9tOJ1Lwb6iIbwg1SKjXJkZYb/SG
/ZSaprEKV2dcRcI2EBq1YjFcIPKB3vbDOe/ZYTkmiito3roPWha54Qfs+fc7XknKkdSDb5O/cU0l
LNWLn+LU8o31BGr0/zeNO399qr5X+22ysEv91ejyBYWO+fYFe6BrokoasAeFd8HCHszI11EypHGL
nSn85x6Iq6xezIyBih6d/uD6/5lhPbuYaq0mANmxLj5wFpndpbvEh/TxtM3KopBBxhTdSPZgHMS6
NlasY1RogkbAsUKugOlhocM82P7q6tGWGkdi11Plt/5Xj8/2AV44b/xg3suJrFovbevrQM0XRbUn
DPppHyvWR1ax8gYm4S4ANVem84ctJldgY/vhtuITR+3cQSwsjORQZC3j7I9e1+Ex2tEiIojWGS/c
1oiKctx4b66kOZ7kgM0zuGr42XtMr+SVScbMfayqrA+rF37Ds0MQA6tzfQIYu0hSa99SHs5GknH7
iveWdeQ9gGRfiGJDTuY2LC1GV8xILh+VQMksgMkO4E+A1Ch6nRgFpj+HWJ6S9rIEpODZRSgtMDHy
NsyRZaYCVHoZ5nWjneYDNizXSktwhulK0ibMMETUxlxw92qkXUxKf6rH91TwPpZFw+2og9e/HPon
dMV4ttckTzaDXzAg2XbRVKO/Ww+vjCCtaJndK0ibK0VQRbl5QGj+VtSmO3bS9r2D3OvtylD7FEWT
+CSRla7ZDj0d21Ep+TsY5nYYrmdOaBjXXoHjV3OaJqCnTK+6XN3vBlmcWw9x0lGMjpjQVaLb+gXc
cG9ZOvnMEfZKVkgzBZ6pwuEoPvmlek3Ifg9nTnRaNnKu1LLur6IFc093Y+rdLU0VlRDo+aGcg5QS
hEnEmSwjkYANS1gsf2fR87KJGYJfdcCbIVAZLOiUu7+5XF6mfyRNwb7NxraVBLB+ex8m81fiMOWZ
DeSzpCXSp9RNAPa3x5Hu7pqy8li+q+YxnXLKlnOfsCW1THl5J+B8QB6z7QMg6nnJCPVCnM5yYJ4k
TIl4p2Odrr3gzOH5Y/PqF5ieEGYxAUwpeLvqPTtcCQM068ANA/XAIeZgLZO9NqvegZ2KDnB9kGhp
gezrhzTVDCS+GF/R9YFxDSsRaAzvglYUdj29+2EAZdbgoF6vYzk27Su4yl/k71CoWcI0/tOHSvm9
3ivoqFKqCd+xpUg77M7d7THGfT/TxGnodstDHfYT6F/JrvG6eBbhD4wXvcquMV7DlF9oP+FLJ0Z9
cqVbkbpal5w7Aw2MhYZCyP74DV79xJPMVsr9gBN0gSZPvpLtwGJv4LPp5KyhRcNf45XZWFwIW3my
a1QP9Z/z6+E+ukt6rd/yo1jrd5KmsPn55c+2jJ3RcTggCdywoYjK4dKmtjOCEPFZ+wbA8zS+SE4i
xavUCngSZxta2Q0fqqWTSqF2UqqkaEpTTrhpSOHICm71sWYeCa34tnkkuDPc+cmY1FvpJA/+A8MS
8NgvZPK81iMxoIyTJXKD7isZKq/L2uhTHNM9xQuqpqCHv03Jll+HlKMNPzVBplJVmWQAYSwSEKGS
60iHT8pnN5gGpndkATJZXb9PBbLJiCRGoNRNETjXZ5Zrs3aseB0buFWxeS+xFzM5de+O0xUg50b2
qSfFPbHykUP737gbTheupqKShrCiSTe9kniChYk8Pbi8Rr5YUYAfaRJL3yWA/8A+zf/aquhDuVnW
JfdM5HMuJ14iDYLuuH0f94x0MUGWlq5/bUcx+hgSsLiSS6mIPbfIgh0NbFaF+hwUxps23088Z0QH
L10HgIXUeGjbSQ6j1tFzG8dCXy1LhkUeZioQfRCB0zZgRJx5WTcUlClXXk2bgm2HF5emAqZNctmC
yX4oZf7K6AE95bgWPqpR3pO0N6hrsuhrXVI9obCgUhEDQ/OGM+NiTbfe7xfuggwAqIf0mWQEICNN
UyLBK+z9Pq3AXwtbF13MOiH5aTij6+ZDJI+dh2mInzPiZcVgVy+CQCemJlsYpX3Kh/EqR1WXdqXi
4juO4qolzrz1BH5F+hWJXm5wgJTWTkZ/EfmPhwhjs/n8XE2O6ecbE1lLB8qERytMuLVaSbhhokCj
qjh5LiFYSa6pbxKAVn+yaOJ7RTo5SS8Ts9T1NLZLxLTT+bgStqIv9RevUyMaHRg037hRLKNhKV2P
PVjFaW+4FhnHZzuHxnTbjjZvXcfpStt/Em8yTzUu7nIW9a7dzW7aVcTMMZGa9VnRUjg6ZufMeJrM
BrC5cty8rToYQ0QwuKq4LkHjl26uOn/dzEI7CQvCVUhtplXIBIIizxsBXhi9IzhrJkfN7nZ2yHQo
DCTCIUTRAGKLbSLBW9E4PDsL5HD7Kc5E5V+wO5sR46jCac7UrbdYAdZxctGLqxG7GLZMB9JW6sN/
Pubd/ymqy86jEVJX0oHQwW0YyLsuBWhp4kpMZb6QLxAFMNa9RjkrTXwmcqQJ47CWcsPnlUQ2SzhY
JL6vZzW5vsJAAyFUPJOqj61lEhgRbqc9EaBkdTj9HKjLKviPi3TyNIpNQobDeFaJp2v/PmJC7Sm+
3t1ZU7wdgJ6Z64dKDvUsQtwSaUc2xH1jM9KpYGn5beVbH6vaV477+7+/5InIcfxYOvjARytOH8u6
cLY0UNCOqaq3eKGHaswvUX+cTkO1fXPxcJiZLsNfjeKBBxq/CwVkQF1hhn0oNRBi9m0QW5oiCIdK
2f7ESGd8630ZXcNmD4cJOfm4+oJQmnzZl9DqZZXZfQ+mx1Ayw9Qck+lTsXQb4e+k54s+QjJDalqM
EhygSlcV8pLn05dijtwSD43+Tx/gFrTvybPz2pAE03YIgGudsnvUVJ5Rr9/PnP//I9KqPPbbUcPC
adzsPX0SNhpHnttkKU1WeFnj86fiJrYuJNlyBlVR1KQ/7k5FuPZ9FRfUySDBhK2OgOv/Zg/hHZCe
TFZ2M+NO1unaJJkchWDPL9E1F6hp8t3sBiyeStGsv/7uuG93uSq9cVSKOUGOCK8lNOKyyzZpgLT2
R1/g3RXVcS6wmP+B+smO46tJCXvE6vi6/XdOa4k4PdDejtdXjl4aWWR/IYoRVGn3YqDcXo8ZyoiQ
FGSc5fyAoOmYBSMQA+wrQ0WKcI7/Z8t81A2F0GqDvyd4/DEb89oPnP78s4ICKtm9mbtcY/na7bsc
LVBQpFb61aLvHwATpUqJmbuzLOj0pDkstCf082TYn3+XSD4w1tLPbcC3cy3O9U2IPXMn3mWzqe/C
Y1cVeZaY/03bqUezAn5xtEwcSIGeEPqy5GCorVervr61pVo3ueMkbesf0Yns8qhsZDWZHIHtpMQ3
JHQklhLZyzLNisYJma9WLXQi36YKfQsidiw+X8dD29VD9+sfAEp72FG1dP4AMQNiNs77nVGwyhIn
raIfCbxz8kG2ZCNhIX3sUDxibY0Qz1aRBr9D2ucpXRz71HMAuWULIfcrvE6re/6+75ifNqemchZY
/l2jJESVja8lbNKLC+UMzLO1LJLU/wc5bFiaN9OLeKXut0TUcigVufmwur/nmQvUD4qOMDyGm3cA
Ucwp3MKqlTKp7PsR1vjZDJjj9llc9C71p2RNQTm0/MA8aCDI8FT5tPdTiVsF4f9+FnKKMEaSJINB
RmwaUqwJxBMqdbWcGWWb7bqvJME6Wth/a1wKjMiySoUZRqfbwckfF+IIwebDVKg7Jo37LFd3CAv4
5n2Ulqmr5Gv3t6jIgSjWM+k5Gx1z759NYzCJhHcQynddgmoX0LIRAqG2sLVKiJowsfQrnpSJXQfY
ATa8AIlb387A3pW6vEv3JWhMG1h35IzMa37FhDjgWA+DjBBi0PqrnN2l/lsNt1PtKNa+a53kJrjm
vK7GuzSEpU/cV2hY++xBhIAXxKKq2Mgxq8k22xmPspPon0Y+7GxkYnKc+AHftJcNWWhgwkqzvgUN
Z39ahzmyP2ZU+LVkWib+ChnSLIOqOb1tdOYnnEvIwcPNWkvTOpQntvQKtJKfGXuVPZr7rYyWX6N1
rTKBGMP32iWWUjjbnudXLDXlt7eNfrTjRabSMAbY1IANTrQyKg7N2NBVIeg6xXCyS3eiQnLwXOF/
7LJusekup8CAbXBbXcdQirxtsgJslGRCK865Dez3UYEbWgEwstcNT3IvvNteQAFjc3UKtqEKmP/A
GdhbMKRFOo+t8eUy0WwpGcwOuUlcGR+X7APu18b7f+84fQx4jf/jnMgPacsfZZ1unqgWCcvy8484
aKVJFwP7E/5HrBbij23HYV8U+RTEGsW873xSnTL0ETNqDCS9Y2dB2YWCyeFbU60fI8/xGnlIa+qh
6B3ArzckhG0A2cOkoeznKa+6bQXoMj3hbmn2zMbzbwQUKFh0CTuMn0AQdeuV8PVlHkPrC9RbQvJ1
gCZ8UdkM0v0kLus+IP+HS5A+Rx4dURo8G7J1KAXuaHnpqTRfXiUb7GTeItM81gViVntOWKei0TxK
sgjyW2gOo0lLnx8srTqfkFmmm+75F/ITezTUZHbQFOP1BHqUWBMx0lEdOVxbER/EtFAvIZBi17wc
MerJl1mo1PKE/pNd6PZIh07X9kuGzL+GculxV6mJ7LtA18vRJUVYndKD+R/ioY948WtCN2uR+aFz
VglJ5PnpgB8HhKPC6PvqgisJ0MUpqJ/xlXGrhFjzyP2L5kb98jDAmgiJ1V1hHxQWS4jKmUPouAXW
IKikA1TPmstTjxo1UWrGu5Nil1v0/GtTA885pL286m5UhN1UN7ZHc6sq3hOf6stBWI+VSGraBQ8n
jQpT32Rcy4FV+fxPWxjNws/JtXjnxD2Vda0oWZ8e++c1LTjBkvexijQBvE4pii3klKbRZ4K1WR2B
ySGxY2AMIorWOODV1ektJeHE6+eGhH0NmKvQIOzKdeniiDKxOmmZM13xq5etmFVIQeF/ivQdkEeL
qeGIi/dzdZcP/u5H1dgjEd1zlHOP5wF8J5gFTka2U6XTNSs1KiL/HFOttYKb5WK5nagxVtbs7IHA
z1Vorg1U131Vff+asnrwl0ycPb7o+yZVA8X37HwzyiHJ1OZxw2I0KrcypZzoQTDgPS3QvTKhNixZ
psU0zFSJS2i3a7jGhjqUwLxLcLo4+UEfS3guCyCWIwbUFwcbILm+0z/rl9Jhrn/dmqtEWT9Samb7
jN9/vuxg/j5zaInQqiFoOi+Od2Eond5hvRJ6xC5F+ykINiaJeOc2DrJ0mOFgvRY5Qsyx8TVYDJzg
4/TwCONxnGZz1/yd/tV6UHP/Ge5lXQV6/mDh+p9iABYv6S0VWTxFsGsUC9h/IJaBgYRHXJWAobfU
Kox1H3e1MirvXzFdKdpK4TczTxb5/WuahcBE1wgMBl4nSvyanRAO+yTTV3jK6dJe69Squ3ineGXM
tYnfmvPRUi6CCwtXHqr13eu1GmLQ5c7YrZz9+rIvAhERSUPGb39M0KJXgO5ZxGUv0JogpT62bLKd
MJEvVIQSuPGlxnfmffMRX0bzjZncHFRVsUN5GMcAMIGIRxxUJ3WdP9ckmn6G4fsK7Kk/Tz6Eiixg
zmafmBjivHDjMYmNSMV1oWTC7x8VNEbdV4zMTWa4y7eZeU96KjTVHys9Krm2tZDa+35y5yTVm3PD
2cZG5CrRwaWX8iHaTKOxHLtttmblxD0av8bSInHX59R5+LrDJ2rmzWwOw/GPlsy3GHMVb/rsnF0Z
zFCigb+QRuFSGeqB13F93idIE78rtJEUP+5+/lXG70+nC8Mq9v8oseVZKkDePrkYdFUxF6/GAlem
ZwMNqJnvXzbjuPaGkjsX0AN8G4PHtIsWtK2UsXcdEn3lH5UmYRz0qNeaRdXNPAEhl65hMV5kHnfT
uFO6iV0+y3+zVAr2HAlKfa+RWlnIe8HI6P49F6LIk6AuWjZXm/bwNUeYZqOHNOgIvWIQtEC22LGs
SDLg7QsmJsC41sSM33+kx8xPQoorJUeg53UyRUbKmkTdvs3eyxMOp2tIaWR7itZykiwQ2/CoTumy
3lCsLLjcpkIKI3efihtHYagaKKVW5QJwO49Zczq4hgyyqHWt7oZbyvxL73eyegtyHtCufjj1jfva
qPjZdzAbgjMQjRPYjetoP9sUF9yrHcoExlJSOJINRPDw16C9nJo6qddMP8L69PwZywugeYCY1hmz
IofEpZ+sAFkIKCyJiYiJWOoWu8+CDM/iBwUNsHhqwjOlZIIY+Za1HP68ghr8WPoLu9y8nyxwRogW
CVPqsx52pMSn2ODfpcD5HPGOD8h+lXAj/IKtai7y58Bvbet74seiafwRRcA+KhOCrOI3ri/eAV1C
QHKG4nS6OGOWJ2+GA+0Xoy0ZIaVDTOHyFs3FYf7cV2/B7I1nYz2Hwm6H0dFBv/XOaOW/+oxez/S9
nKThaFCg1zONAywttwUZbTkpPwS+pGTdvN+xLnodOqqzbu2OeUAvjWPOF/oX6KfkZPOydSRsL2+O
m5m6B6YA/YY17MnPWaG89pli1phEBM1H+x+qZ9wrsmwe0RpInv9lf1OiTQoVIHzwoUlJCjTpRuPF
T3BmBbO2tjphlRLNa4DgtSEA4wVXe3NueTEbAjRqZzstFgI+17QxdCeL7DoYUCNFncLAHxNJ5iif
sXYNVQopH+wDgvJwRocRGdtz81BHPxbbwHa0c7XzlD3es8mEKnZTn8Z7kLRyNdKMa3gI4fe9WHvS
z5E7A9aUOsAavwHOw9BUU/Ozzs75nnR6k/FaMGByves2PsTSpmRf90l33l9tVK73ArJmcVK/i++6
JJyr5jYuDCBDapc4ysIoIbuTgsIjmX2wNI43fCbKKRDHJxprmNxJ+kNpWkeeDUqXtAL1fBjiZm32
fYBwVB8s7n5TeoX2NWjMAraeZFmBgrU1t2Z+zHUD6qXwWBmW7y1O/I4b/rVAYtqQ0ZsjpFEC7Sfn
H2JoAP0YI0QNuxACdZf+dP0BAwSQlXzPlInPEOce2nRKHdU3UHhgUx8CmT4DAGAhrv20ZCHZBwFl
5rmIaUr49OJhCURY2LyLT/+e1UixaOzF7Gi7nf/HjpJp1Fr/obuD+c49VHcBifF+zw0t87VIWtd/
p/XWyA9YAQ3yAmLaxMydLD6ZuHtk6jMASEiZBlr4+faiC06zGmn9l3mqMGFXBwmHAWS8xoBOE78D
P4PhjNrO9IaHtVWnHW5y0ixmI7B9WdK/TdRsIEDTPf8Q5JiCl5ZEjLnILL8y/BVqpEtGN+qIMsVp
Qwf13cQhTulIO74eRuYX0D8wUcJPiv5iv53gVb4PL+hdRKkp758/YW6ZcN83WRH3qUdWdZ8XOtOY
ubUha+SHrB/UybENQw9Um9lC7B5orqD6BkVcEAG7lFDjIjRE494T7TJADkYqKPN/au4xRCFu4Ca7
9LumQaj5SxYk+ZF6jfEMML490Oei99/t2LR7Mf1djIDwWo5rPjhB1x0oZJ3IspLf3oFF0Cf6NjVl
7U8gLHcMDFVo8VZ5BizMN1MNppu+RsR5/jtFuc67VfP5+ltdjR2LXJzXvA7UaMpCBqKTaFiQnNha
hW3uPoN2jv+bOsf/MWqcTt8HjIbAZgJ7nM8xuH9+LQ0dCzN0b0QhPd14CV1FHssOQzXVd0KoZlFq
Xth9CaQV4qJQoxXwjew6j3pJmK9JqDmtjFXkaoyaeozLhH3RGYpU6ecc1CnBophmjbOobVW7dvbX
hZ2EFEp0Dye4wQEPaTUIz5Q5KGntn5OLkO8JuXr9NY7u7TUV2OtUVLsF0AAbfjq0uq390aefQW/c
2nYY5YCWux2N1c9/OCRdyYn4IDPWI8lZcsOin7kmuZOaSNwJ3zQPuh10VGk9T1qRRHN1ZOqSLQ/q
tyx0Qo6A/GBptg05AkCyeZa4LYj4s/rVt3yOIEdkX2SQ/QJZe8qM+3yfkG4t2hvlXeTTr16En0LF
tRhapl0gCpYAWx1pgu7p1iKN9nrP4q2KGLmQVmmBjTOrPbac20zgOMTeTrVWUs8OnZQfFl1exPv3
NOqC9usVt62VUMZszydH50y8klCPm03p/pbwN7rGpLAq4vJBFLKmd6cY48gciLouJN14kpTqxIu+
ABVwIewcPTRs8nAlpPP193YuAjKiJb6YzjCxcz6hQNMqYF1didweLi+zJH7WhvqmLYQbeT1BMjZh
2PHjPQajzoEljxcKUhdE3UB6gSzyXovOEtWJTA5TggTBP+6FjdXitYI1992KI1ar4p+bDJOBp0mD
EgjaqyYUTUBkwEiSTDJ32TcfzwSOfbr5KbAvYWSTlwLxXxf+c5/Wkv0pUMXaFsr+8oU7TgUtOWlG
a+DmxTvyRsSIa8T+voxHT9SlIbMDvQj0R9b/p6rikfM0G11OKcGuDwOsXFVr7EwEaMyC4KuNFokn
szioHCcneCoxVy3+qMAXN2NZHL4VbPwP4WmNqSr2483kLL93I7drgeEG8ZO5Vh+DUvZrfNgdBjxM
v0sBV5pOpZR5LVJw8b6I8NfgXjHnoarV8MUm2JFO8WsvKq2RXyqc2q6ajUh77XTawzuwK05KGwpN
fUKZyFzzVC/TEiBO6FmrpHvTrUAO4geZrQyG7XAvTapJphpBJmYDOg1lwaE5dhBbamK/px9g699w
jaKhzgbqQKqPGc8QNbBiymf8FqX50liRHK4mRvYHn5mXQJg5NNfPoGXSLabo1MYcMJl0FDXim+Xx
fK6z1rAAUyxLDuP341bvbWU52i2q25TCimljRX+sOHU8dxGr/ZWlSY4fzuWpnjq/Fh149XMOv2wc
bkHrjWDI0ci2Y9+ys5qCo9Y/ihXpT1mlP0r2IITEuAAYiygRCGwzPRAgcF9MzpnXklaD+ClMh2ue
3LNgxZrbc5BLXNjlLt/BFq53+yqnwNYB+iN6bqMS3DRO+lhdeANB9QUoNFZipTQ/h1eQa30pDe/H
T2ecZeRbGOFJtBV+bfHxUJsNgcHEGqwKQpTkj9fJWzlu7NblMN9yAlJqd2yTPOqikZYI4BwdfakV
eCAO/zdqo/ajlvAQBcFe9GiJK/VYP8069kuvmokfJisRgtJsq5LH6bVHRn9MeSWk0nskOwWS0XTi
HM8qF5G2FY2IZywd6uXtQdrJNvcmUyiwgB4EOQFI6sQP/N0BGzjmZu0vbcGjgKaeK+0sIYCzrIT6
LxGtwwFFOnYjwoTazrzV5n6/4ll+Pluo02L9YGPerpWr2S/wGbsVt0QrxLNIsgSMXpM0mgNdd0IM
O+BcoQR7MZ9/vKbnNqF4TYSl9gSrm5PyU0f6m7lwXuVt+YkztqQQefIa7DUtPv59M/dedBdXRz/2
9CLqwfH8G09bf+ZeF9ngnhTaapQ4y1o09XqTkYD3RUiYCfVitCpiSZrupDwjf1ukf/jEjhsDfKy2
1no1clU+7UrR83RR6m25PQj80+Q/dhWte8r2p533F1TPvvS2JN+GObxniV+CnApejBJ0w9KFIUFj
5mMbLHX9fbrz9jlwQ57y8u9I0E1mK+5rIFymqGcocMGqsk7tbajMlBYwo4nSkObxaYrgkjnIouMz
NFntJ0SUoUUHWeLaLvisJQMqCVAXkf/4hRMh3g1OmOO+iSwbG6KI0hgXDMe8QXPMGXoavc+iz6TS
m2PdShE4SzZszjcz8LqgJ+LyBTRF0SCsueyCqU6OZJsgDauG/iKhDL2GF2uK9blv7alaH3cWx4r1
dDOLPpKtwWjQF+9h2qXbyGKGEXSTJpigsfWTazxvIFum8jEM5gOUA14+jbbyIYhvmKRXCOzPE29i
iZi9fEpuHpP2xbTpOuP4TBxNbvPXNy/Z7UNfz3f9CUArzXz8phfJBzOjX1RtOfp3xhw/s/+iwtGG
BWqOmtn2sydDfTYNgopPGkbNNm7z7Q1Z7+4+KLuCQ+wACk45uFzB8vbgeigVYWnz1gyY999e6fHd
d6aGyL3yGJqakwZv6P5qnZDAhh+eat7azlVGx2bHa19GETodxEOxKaaFLm/2NvhrWPbSGawPGMaN
MgQ0Amg1FST/OKm6GIpHMeHMFXbdAkUZnJMQfF68pHUstC9ghRdvYjr8igLoFHVreiySzMmz7f6V
+iXzgFdy8pqkbx+zK5Bm4BuaxaOA41ImnSIbQUr+Aaf138WzvUAkHz29V59VyHOrlkYVTyR0whHc
/r5FMKUPbBv5381+xhKa+V7/lWkDsLDilAlMobxaYmIz534B60Vpl+SYVFPHbapVcRekHb2Noqxl
Ct2B9aCnAMRqZ260Sp8nccSIPqMI5Nh8kwszmAD/9usBuzBhBcd+Su9wONcDtA6uAbnj7tDCDYw0
aYwli0r6s1DGOF9nwNuplk/PW+CzIgKBIBNN17IYZi/Q/5/yW5Xjxdag/zHyj7zPER2hcpimeYJZ
LTjFDVnbAOx71eDkWBkxT3+dOIE7WqIcB/XJadr1YIh6tpJlNdXTbyoU5HYWgyWPkAyAlBQ/Cd0E
b3JgPZ648Ja+den3M7/PU1HYLSStWrolvfVejNPHrgF/RM++oHK2DAf8uaivbVPkCb9Ox1BSOKu1
CD/W41QiC4DZoudcRvlGwsmIxLoNWAt15bfQSSucKM8SVwU/hw0qRqe/aES8Wmr5X3H4x5I720b6
4qP78Uss79vv5GTDuOfjnoY220OM+LBNH4G1pohTQGDTyTX5BDqH6EClVgQHRx+F9GB8ZQTLyYr8
/h7PszR6zLC8kuoA511u9wKvULqHxDd1TAPHkNSWW3TVvT+5xQZ5QjMeQiPUkrBVKtwRRMedSbAi
HW+Ocr64hBIFyT+rq06RMT+J86AC7N3JN9jsR3qu0oS1DF4d/YmoHcUfMwv8M0ShG8Z1Rw2je5U4
SvXlJY3zG8ZK1pVIkNB1wIJH9PBl8EgdhUG0kvg7WS8XhmwCSVoyPuR+lSfFRhWDFZ7jMSdYwci9
sQHLYri43lcT0vgioHHPCOOZ2InQHx+NiJWiIvQdMhQ/1Q3Q8wBrmwDZfvGlVxWOnuBQPZfi0f+w
9TESwW8wTrMei9JGEPg2nmvUal0bXlEK7Xc3Md+bHU/lq/XHJFTT1BTHwA02DBlRC2JKCsR1R2Kj
/1xilNe7Ami7Y8F8AvGScEvUl6SPlhAtYsBtKOaF4ryi8HuXUcgD1x3nISh27HVI0PFbxEt3o++O
IuY1iQl9J4V3YxRybcRhtIAFQyAQ2FjHcxpJOlxMiWM9vk39GIur6kqVE1zlu3hTKoGAp/xG/z1I
0CFyegD3GjfvuDd+jfK52ek9hSLPnaAhxNSpBybiSQ//y5c6S8wa98u4sgfwikF6lBDN1XyIi1VH
q1E8ckTj57Sfm4mywW9nldA3IiH+5EDJfbZ7ACRFR6ey/RDAwX55umtdIPoZ8VNJvkRvKuixfvV+
JOK3c4TIx2fEk4Ae0YuCg6ymzpDe3y4SWV0qDRaqNY88iERJjHoe1MJcNpznY3xfZwamNdm34CTW
KE6leqHk6OI//5areJK2dUdA/AO2XtHrYBnqS/eXChhnFxGNzJKFdfAbA+jteO05cur24MdDTGjx
DMf37j4ldX9z2AE5sDwgKzhMd/ZEn93UCb4tCSLVqdEYrSr53titxnNcseju413TrR4UW3cuwjwI
7OPrWq+nMwugl4Knhse/rLhMGw0Ok1qOqjLioE6yVYbo4jlNQKI4asi3O+X5wsbQTlZDba6HTD7g
+5We6qIgIINa9BG0S0ybeo1DzLyzKGnK7ZF/tj4GD9GdA++WXX9BBlK+pLWQ+UCM3IuyKlYMONPv
J+u7KI+Ah23BQhCc8z4w/JNTl0ei2IP2fkvXzixsXxd+j64TAyzxpimKyK6f12ouQ3F+Zs0v2L5O
zpzoJIZXcTet5VGYzRjBy7l0OXPaFPWkLh2FmkvpXUnid1ks/JQEtRHBhBXsGg08ZkGKBC62yTMv
V/Ltpr0vYptadgTZssoSXbFKBk8UM2+BM+DeEhqFVUOnpgwXKoRWEjA9DLQj2C8DRYVuwX4cLf+j
Kj0VHPuH3Z+GyKrftw4464KR48LySJ3hj8K9e0wuz63rn00yRnVaAZORzPCOGd8AaMeifmV724Zm
mudstc6nvoJerrmnONTdUnmeyftpHpi/eJACUMp7Gt5dWjnxD4TyHtMEf2mD2QPuxRfGd0PRNx7d
g58VlOHeJ/1PSICkE6dZYOrnhhFKmQMSmCB8PFV6/9HfcGBLVIS6EQsEtnw14P7SuviezrwW0b1G
RUak2YcqUnrn6n6aHPZkvDfki/vxsYA3UnOxDoZxLzpiPVeACRt7USz/Mg9yyXTxVgLDji23xm+R
BhPSjFgw2PKMjspQVgWh7vIVnnKS1AFRqZMVIrHsfdZy1WCOb8OWn0dG5Yr7IaeFsUJAaCWITJJk
EeUfF/OuhtU3klGBg4FW+R+M5lwdAPzeB5a3YGdGPpVIEcNIH73GgMTmj4plS3zMQlTgAcFYgRXw
kZPCht33l9WZgbW5ecqg/fRHe3VDAT6imJ1vwvbbFFlygd+PamfUyYYMdumxyTkQyCfh9HUt+rMW
G24KUHHsTO99b8Q7TTaSqCxDbSLv1lDbGwxMquOahsBFvkGJbmUAReAFI/Aj1ac46m6CvrU8atVh
9mW+SX1AEfrnVu2UIRlhdzYpQDKWHCLFxPIDAHT0QpPKZ/jjJz0n455Qm1/UJaSflgHIlkBGw3FI
62WzyvuVK2aGYPYyHXS6c/BGpvjELdhwr535hJsAZDnFcKmk4Mx8/xSAtXnDXQjKcgjkT1ICEozq
AaNiPJiWIoQ95GXc9QwRQ+CXri5QAY/dyT7w8xsNdqTvs+gSaDo9oNM3O3jM+yU419pvVnXVYg+i
dnR0sK6wvWrijue5ZJ2rzDxRidO28tuJv7lmrpGNKSnV2MmkSXUcJQMb2QBS+7S+F6zM2/ofdcTZ
zNvbsxfjd7lzsO3dz7CQVVL/5roMcJ33sbHK5EbMds3V2k5uQ0UarWXmNZrKHNQNVHCHBj3754RU
+7i35L+pVWRR5746N76fzWX1FAVa+L3h/eYXM0sdzXOZP+AEr0OH48NpCCRMrQzQ+gCJaO8MUq61
T3E/3GWClzl+U6vIfZWyLsBXhRMxVqt2AhaiMqUUunwBOl1EAoUwssjLRR3QddORdc0VBnCcJMQV
teLITAhu6RlTSj4FMkkPjPa98DrpySakM99mlwxgmtZuIvpJXy78C378ymEXOtY4My0BEDG/EVEL
nRes8q3X0xiX2/cp/glkwpsHwCmNywPwjsAVsQjBcxJ1A+AwF7y9v0xS45h/4NfnO40CbTwP1mLf
vH8DVFyIHVcibrGM6YGfQnQLWnby/ccVakbhFvdU+XWFqi8mb0VuuOZgKVC6nodgXLx4gaPPyRl4
Pm4Acmi+lNak882Xq92q8hdGnZG0Czxlz8YNiT/W3jzaf6oLQ5oL2j2ZmB2ty0PFoBe5E2Roowc4
gEq8LSgx49M6OlxS/GppD29d+yQ8cFT9HRyVYgHbaZ9gIyPjsWLzH1A6jZLcmC2ccpnnUriFeBTK
KW+/xvovc7m6hjS5ui8Hpew1NwISdcfCtYHsRMge/0ghxOIv2rb2pFgVbOAB69pC8Y8dg2a/TX2q
bFffdtPfctJ3FcLIv7s76iPuhXKDVuGEqwlxv774wSchgyWswvaQXCdO1UQI+urMEokvUwOMsON/
Mju3qxfOVWECyoMg8LfxOYAAebPmJje8x6k3VQduKpzHuxwqjsA7dg4ZhV9uThRtr7JhWctvpgcP
4t10KE5rBs9jrjkPnPek0RjaXDv2sZw14f8RzYYkM+32xZl9l/I0fZFpHLMafR90kT0hzFI9bpdx
0TNmUXcJrq4c36a9ugcLR+Hu8Mxgw9wZp6IWhL81lXEL7g0ztgUFy9gHMBo25prFx6GIcPsepJ2/
PrGDjHaQCsCl8pJpIS4vtBPAdZQfnm8OETUH8qPp6B3aXky2HoS3VbClmvdT8Ec5i5rc9EjDkyNt
uadi7w2kUfhzGb+63ZFGFpFJSVQeemClf8LJlGEaKkJACTCX85N2mdcpSrO61TP0hDPeYFG9YN8a
i5y0j+BW8tqJuNHcLTZiVmbpIHizELdZ2lJ/6rtWNL7kq87PC0tCTYwgiCYU4SkTYz5yBYzdN9+7
OcLXJvXCIze5q9NVxkz392Sd3SZCZMnIvL0YjeHsdUwK8Wr/f8QoBLafKbvf37V9fr8b7koJAr7t
5yOkw6LyShMaDjcVfr2KWkVGeewMntKtq27GKvebq1iM2poe9N5yf3ZeHvADO4UWoCta2zy8L+/C
CmCiKmsCezd2bquin1EpPYXIODqIKwyxHLmHBS+lhzWGzRuG1xWKkZBi6cVuKrOd9MjEUwc6mIAn
uX8a5aNXVyFivfVM2iBIdkhLGILHH5iDDUQF0D4xb5iTrErppe0Cm53cbz7NghG4GSXK+3Z1t7i/
d+rnYIpND+ezsgEF7to/+s/OJ+mKvo52HMlt1LRd4WBNPgYKBrz7jzX/3uQVAvsaEiYbfxhVG68J
WTb+Oyzz00xuAx5R8qG9DUtSsCDy9mORnLfmRRzyUIkqFu7s5QWtmOv4TnOKWATV6WvBYtje7+Bo
81Pz2lq0rDIX+k9CyDF6S9oj1y95laoxL1Ukli5I7dfsNV5jKnpbnV0Eb47L0AVbI+1LBOlf0DQN
pUZ1nAy3/MdZXuHDFfkseztk8sYybPbEKICkL6i2RBrn6QhPPXJdmyCabgDnMxgU196maOYGWCcV
wcuDI+PyUBFItxJ8B4VtBHko0QmfrDHR84fNZbf79Zdf47qhfNBFZ2gCB5yPa8UgACli4wSjUNRw
VovctjXO/3qd4qLnBoz8Ao4twJagTvfEM5Kqf/VpRL5/4WiIfyFDEuGDXhReHDMb11nhvI2itWHU
SVnMtsl+aIJxQyjdaPjbMJaI3ap9fkr9XOMadZdkHwtRBndaW1J+PNoM5IBKxh0w8KQJrEDgbFpI
jWZPAWeZoUotdWiXOkYi9ltgmBFXJeQWL2B6eHM5vG80IaSGtNg+KRhoD0Ytl/McAsccOr3kgCvy
TCBVXoclwbHzaVTUBj4n40fc+jrejj0BJdFRMdubxsPejGIwZt0eftsnPZ3p4LCZPHBglatjzCBG
D9enzKzj1NWjkBAj4PY/ch99YVVIzZKqrDhfKflqqMJ2xrHpBPW0kHSuVFUpHcZo2iv6XYxgwHSF
e+R4IOUCcoTYBgJ8fejszcVJ8dBajUvMvA8ClFryO3Ce0XnqDyVx2WibaoETWAWVPrTuSXFZ1+46
9cEkjP5941pSfoArdB0ORhzBhxiF9PRcJhTNcw//doIf+yil3XsTJDcPjI6R0LSOOYQvlzzIWm9R
Yyy66EIxsr3bwEavwYk0GWBe9NUOm4n83w50rIMiMTL7qEXJGi24y1su11coxWQME5wrXjPqvytE
SqW4QZXttGnGXHSL6IVsgNH7Lfk1LLAclE0yyn1uv+b2cy3SRtmfkQfMSAaJtsEUQcsMrCTRiFb2
F4wHPKPG/15CkJl2ddnRxT505ZGZz1YrLWP1Ag8QbzUj4je48BUaoV5C3m5M/M2YnFqiqfu6SRpE
pf6trktoCOwcP9iSF20PwInpPMfFyGCfarumacyVMYLd5xdJqjhk519ImjRMiRfgZWpSJqiN8BXK
Hh2r5o9l744hOI4bYnoX1Seg/opUPMMA/itcx8Q6+xmAjPgC6PxOfmS4DtUTxJ8oxbrzMQdRi5Dm
YA88fkKx047gdn15Ra4sj4l22UT08DGbSmLISorNbgefp+/xHfZpAQn0S0vIdhtfXxzsPOUrT4md
gUhLdTpwV/XFTQ0xbyA5eNWJOpW3nH5Z4P3uEwO5TACYiLJ8kJSYDm964+3qn/EGzukF4hWhVdy5
VHNOo7mknsfAcu+MXn4tJBnHAzst01JHFThL28cKQQu7HGnbNvV8GcyHwjhVLdmdFX/KAiANC2hg
pJuPOlqpEvAhigqbrAum0hbdZaSz8CJzUzSbQBQRdpoqcEdg9uOxB9V1NL9fPO3jX4hbrcJeaGOi
C4PXouZfFG1l6CpjiJKrBOjPik8wjPaWeJKaI6FtGF4TJQJ8gW5SVLGxX/uYzOzbF/1s7pIrFsGu
Idb+GEdyZ71jjg7+ge30ogy/yBA4ULqHXqZ0NKzxksnXDPyDx0lkG0iSgmumKV9zVImQed7/uz3R
t0Iv8X0sitjPEiv+NtD832h3/Q9k5WQRNyY894iYOG0ZI5Az32/eZAS+Ucebx933xhY7rD6B74mK
7LJqxE2yZRoR01tegX8U/qeTnAiaEu8LfLWwQCr2YyTmGffSuqFfmar1N8X/g8ENEdxPMTuGi6wF
dhwUxWTx8/sbrl4EnNCtcjs7M4NrPq0Ceo1jISWonlmZmtEcP3SdmVhnDSBpX0GpUOxfYpWGb7hX
MKpM9796g84hgjsle190WnQo27G4ySNJtq40UWyo/Wfi6bbVe1aP+pI+H3gk35yOfIF/te4/47mY
ecNwaZ3NZSvYHpZ1e5RvBflGM9z5DV+S8xUpMovmeiQCtx75uu/wXFnSiENTgC+GTWTgmAO4J7tT
VR3NDejIBhQTeTf5yQjafT1oWFyBqgJkuBcVKMbCC5RE/lznXTLmQRn6z1r/Ffj+5vNmBOt3bIPQ
GJleKYXGXzqHpouY3tCkTygrdxDYwU9Q/SR5S+y/AACuwqv/ycK1IG5eGVXzOfHd8xBpmFQZPsP7
+WiVuw5qrBbXkPgID3NOif1SSUH46mqHvSiF6oa+bSF4hclDMln+c35mNAseJhyEvQNCA4ZDw0fK
5/36aY7Iq05i1dBKYnm6jbTboLelzfZJZx4fElvryNqIP5kqN4k1anZpsRt5hMR3Ff1kHL48wxKY
xUJcF4rpJaqRKfacPhhKnbf/4bKnhnDW+HS7KEgsiBjDSjrHwtcC/MEVnNS7ppwFwHaCghZzN2zk
EhaU9uQzLdmUKWUBUpDodhsAoMHjYXnZVJXqD3su3nZw275nh6MmC9M/rEqZNL64ThcFqDI5q/ps
yW6y0zLI6qckRtX0MMNF+iZGqV5Gu/+CgOnOjfpWsivq1FvHOWE5jdlchoGipEyLDbnvCrNru9m4
HGCAnld5zikt9Lji8fxGsfU72zVUGUTPXqKY3xrOpBiCRAcOaetB2gochXErqsu33Llu2afHXcpR
7WKVP71n4do9++0XpwkbIaG690Vkyo3QtdKDfE57QboKLMxAcFvXZWmY8nIKBU+jHEKN4CtwEq7u
ZUa10msRf9g3P04silT8sLSF2LFpOAfyr9kVhzmOsnxmXAvZwkAu2otmy1WESrlZnIDkBXPO0yMK
xelFQWH32v3PVuLUJzyVV6lXMacT8DjNOxYM7F6gUHOxH1GnutxTSTYYYJmAn2r626x2tLIh1Lsu
7KPWyRcmkqHGesbV02U6JjwWv1taboMofkABtH/Iu2T1Lt/dD1V6I6Se+6ub3yMrKFQOUEZByzgJ
QKGUUHJQxuzhwta3abMHTC1LZyHzvCuZbjB17WDuegCcyB7J7FblYVddNPBoMkriUAu05vhFroCl
CMUQuarySUSvJF7/U3pQzfXkGVIOEieVng1kW5owBjxp9e918Cbx1AikcuNbYfMcCOH2SeZQ845Q
8z+uU9k/6wwjQfSJk+Te9e4FgYa1+qS0BKuhUfwbaz2wvcWiwFY4qUkiBDwWleepH7AFudYwB2FF
H+Nk9inieX/qZmNSohNLSSwLiG7Zf47NRBt1ChvOl53yxjUFKmKOpsGYUdv2ZyXrVavhY2mEYaM9
fY9uwKDOp7qZZRITkyIjneEd2CKlJgVZQescCA8lpmRfgpc5VLCW3t3LIIxPSmTupyC6o+5lF2JD
xWr9Xxy/Xcsr4U4XAGpQs2wYRNplB7CSOKGIjG9u4lMBSr35rLNpJuCYeT1VnlRHy1lu+4xQQiKM
OTZYiGf5bakWRygifBM1IqB/12WWcDSeLKOntsvhiTgIjbvJ5yN/EXND1afjXoeR1NuTrBX/a0Mc
dcs5bPmg9ejRphA1kx/7xqd8qcfV4dc5D15jfMs+52/oSkIzqlwuXw7BRdtlAw1ztVQiZYay7J9Q
qLJJVp5moaFu/VvmZb5tiUL6Oc+4BtZXUitctwFNv52VIfIwyoKWDIlba1UAucN3YIZcUFY9DS9e
j3pZ+Ro1cndTh935KBihymeRiMqnyeShxrMjnPmQLQ+usyMoWDJ71mmsKeHC/jlFFWExaUdIVDWw
lcx7fQDpniiv8tS/szhYgrTTuiG4/YNpq3k9PfYtRxNQD0coK1NG/CWjTW0w/Ijwpec56xRi4t2y
gizg6RXHsOyLzMqjl5HZUETsOegsP9D6rnjusr/3QmzwLq9WcQwqxMW2XgfVRzJYhAbIx8WfTsd0
PVNsJ2SFP1VsIVZR5MoblLil3bLwPvhawDktd7O269z9TEt+3ASMe9WWU/5qh7hExe4fQUgylAG/
jk5hZPE+XoqlqssXF4TunSPheDb5SrWy2GB0OWtObi/JCKf5Mw4fFLbbtYMJ5K25lR1c5+nxPh1e
laoFr6bb63z38m8aUZ4eIHv41PuAaM4NrG8ALtA4BsH84k/P2TZIipWcVJ9A0KbeW+zt8c+ndqXh
orNodkPu6KFPp6UkvEfvkSmEzG/xfhiG/SJFbVWlV/ldtk1vtkOmvFeWrMIrUl6DXByp0XbLgx0F
mKE6ZFCcYWMyM/aJQPoZOqMV90QyjQQ9KnqYhabQ1AukuI32qmYMqNb1/0MWaoLyyEO/VuD7FLjO
QoIR3q0S7WyzBnCuBCqnHW4MN673RCZWlmMb3PzB5W9LBW4lmmOJQJpuTVXqGmL9AbYIlbkh3mhq
p/fKc9gQ0KjzXWIhISiq8C1+p6NPwsFMfV2VkoUQz4E8H9hJJDzCufP78s0i73hY9paZT5mRlJWq
QsG8P/CAM08IGqcJ+NfCfiOS7r3NGbe5vTT+AxUZzetuUmj3/FFT6REPsi5CFu1/0JauBPvU7kz/
nU1Llpxl8Cn9/jiIR//JOi80CkWy+au4gooEPFw8jWrZAUsT6MMuFMq06ZR3new4I190Mh1CPCEn
vnE006Bez0pc4Fnf+f0jUWF/Z40xeHxT7d2VT3Ww0pIhdqDy5lVGOmeaU9YP5enlUfBm4MNCNN8K
eRgkHfmincD/EOEV0Cv56cHDtI8NLaNsB4XPPdMXjwix0VldUxMZGRznbwq3JdpsfPaxE0RZqvEN
wrpJPboNlTH2GAsMbD/XWK1VcNmig1asi2WrX+cV6fBbCV1jIhYGD7abzH8AIyuPqmrobDrSq8Ix
2kJEgptC6iw8aqDJOEqtShtgustjZtaw5LhYuOZQAQEE1zNOSiiApwGX8oto5OS89Y8wVP3BdMPQ
JskpE98cR8xmfS/9RlMNsHhN+O7nRcd4ksYtrwXRmtgNy4FbdMMUwcAksBEtl3q+cUpe7b5c0zcJ
987Eld5dEon61eE6feb69kNCrDliaYEZspIo6TNmLc9eqB1Hag3boFJv5M9Afv9khQH8hvfAKdgx
h65tBaZpbJBbVmmMZlJyFfTQKuJRble539GEThnXDlxR1RxBSnbgEUblTIFJPBSeJ+UlnJzRkF6+
I3kItJW2ckqSOaFVl7a6KnFG0K0KzbV0U8cJwlP8OIJNwHCM9Jl12Eksr/NAM9cARBKapoxcGyC9
EqFxgTxwUYzmXqlaW3OuOJYJIPE60bykfOsVAKHYw4N8O/UdhDOfronv1sWISlo5zRowxl1P44oT
EFU10uvpclnTw4F4YblcC79JvbT1GsG6I7jk4hIzKFwVCGQqY1ihGil7iJ2J+AhUem2XmR9KmIaB
qRuI4sCQarldRUyer34ssNZFhalA+tA2AeKn9+TALR6iKOWKfl9IXJSeMzTOtdCIZHkuB46tvRad
0aw5uOR3xkwgCr7bMH0LQegbJFQKwfl+tTbt+TmeYmg4ZEOdk684JQ5L69Er4pmPudCepaLKrYdd
R8M/GRLvgyjRLZDnctAo7JmLU9wblqh4Z/hlibHqBzzcDl3zM0LAMiRWCiTnedU8eAzEjo4N+xuX
4a3MJ6kZ5tCH1srdolR8LQMtfF2MnG2/5dshoQDmROBJZ1gVjy5wlRfCn3OytpyOU6xmMnr3fxXy
GVfyLEcWLa9QLJ9+ENZiJM0xsXM14Fj5CbQifaZIygbc+fyLHCsv7LD7FInfwOv8ON8dJRLW6+SV
Gg0IR6DURSeKXZnLTXlEdoE5Om2luj5PtMp2L9Cbca9BJgsRB+Uu0ztL0NiDpoVJiGCkncQNzysS
AOWupAs3t0RKCmVMXUpq0GKp8zXqOPoh1rqK2al9Yih8YO/SeNW8G2e0DyoJtIbf/uY/FituXGF/
iY/7gs4T+wVDyPBB5WvWjxXmt+SkO2puBqa8neBGSnN1IbiHtGXlBV4BoXyO35pFJNfcoe6lYzPd
7KC3ZtxJtHN125ZYZ/8avcLWuOzWJWFZzHSWl/1tF4gdY6OYX9AfPoOD4TY1J3AoHeUjHmUPgm4G
nbjelkYFQWw/5jPWlRbnrpZbYSSBJ7lGbEadE0FJzdebbYE2Oc+kmuZFnvSCRyXa1NlTXF9vZUOG
/gK28osXfpxkMjp5lVzNCVgSM4YoFDZSqjFnbImNNzB1QT75sGyu6p2/gYhkC4kiZbM2C0XcNcH1
ZjfSoLFAOlDsH5O/qoK+3dB5tu7Q0vTw2gZVNsjUaEW4tvlRqtM+CHuQr3v50FPaSHo2fPq95LXq
F7ZUmSqgd+mWF+3zm8JErBbrLT7FyBAuqf6U1meqEuWIM4/m3S0ubmGTqorhgA2C3Frvr1rotZg2
RDlQAaMImYGAQFBFt9FdpMhwwblo+aGV/x85j68hJRLQRqH7cDgPz85MiiBYmCoS9CQaIbAiYaCN
1tAreglEqvNZAhT2/cokSCeMV7EL3z+Lf8E72kxWkqjOEl3cEwmEoxu52mUG8LeMBoZiq3iWiKhI
7LPpZYhfQLgrs9ejbiZGKKbdfoZN9+8cGXvnHidUP3eZhKk2qPs2iO0VLRf7WAIt8K+rGcmyxiMM
9tIfBFcRqxjJCyKAHTb9iLYTtptnx4rCVq33qIW6VRFMkOrgCD4/kM9BcgDzXM9yBI3nd9as2qMo
DG9Dg/H4j6OxODTUrr4a3yizOQmsR0p6RH/rJR93OxZQH/11WcqzEaARIgkDrwuVinYGK2ssTffh
Wr7705C2kEhjKK7xV6Jv5rRiUam6JvcvzobuKWsE2jfToFv4r4ZOpzL7SinIV2VtwUCJu5ivvQ+q
fRVQCbcGa//U2B9tGdypm83q1wGJrDxCvySJvBcxlAU2BVON/ytJRkQl6KOouZ6ifpKU/hFnw3O8
hyJ46tpZZV9PNNYHbe8tfeQMO3VZQw8/CDSj9RJDJmbNtc0YxkBDKgeVeLHRhu7PWuGVKGbocaqZ
sX7tbsdVb2z8nEgr0GcPb87viNMUJuYHVezMVze/vAHDjSTXnonbOlI0QWo5lwO1LKiYZc2t0zE0
J3G2JIvfUf7jybSdzAznjLAcY33SpkwFQxbhhM/GUamrQvTyx1anSRSUKJ5/yAPd5l5YJITULyBl
2YfhwmSq1kbFPgqHR5qn1dqkEUfywmNX2Lf1Nvmci7QtaKc1Br7W5T/6cBDTrSCfmZUOY/Mof5iY
2TVVtCyaAPLQeG9irQ/vfMPs02mvy1QON31Pj+UF2vcKi5MlY4Bl1qRJ4dzf6KWcbZUZRF9q8esc
Uh4MRe53QO3pUnQ6zwmBzeOAivB8PPMy1TeOwNk/TBSfAVhWt50gS8hrc2ZzxiyzOX9CVN5j/t94
UHSKTKc7u5UrjvjkHmCw7gIz+cJgZtrffQLyYmZ2MH8Q9ipejUXBS0Ri84Re8DovRsE360dYU8J7
RyY9Rjuumtb9i9sgFCSjtoU/V5tYlQ+OSZv25ywk89Q0WDWke/ZXX5/13ng2UOlMIDhxYIA88NNz
uS30Uq2Kp1j09cYx8FsPcCsZAPS6HXWcOEdVJBAHy0hmSWvhgweJEhvvaJi9TubuWqAtFvJILeNW
6gbDdy7424qxR0+NfGD3fCGny/H3CE6xXwz/DZaR7B2IMtWDl2/wjqrnuXLK/fhkeZae3LH1xMX7
Stfau9qwO7l4uDuInWrAsgS6IW3RHJMTgSnIbxsfTXO7A5zCaSVCXIuitjXkwId+RDCj5oyBct/u
de/r3ga7EpDU4lSIBeVPnH2sj3U3fjDegpgYu3OpJpSY+gChTU6O+Ugomw23nktaHes/kgwZSZP3
US3syYtC37bwhwL4K7Q0Po+Qf3d8jbNSexPTDitNn6KXekmLEMVMeP+mG/uKWQ+JDRENXtO22IKO
RrM4hTqjk4iUXW9pASXMXCdcoc+MAbHDktQdjydlOTvPOxMDDyCvMJC6ykOW6zao+mAqhBNOxw1t
r1jrwdVQumiNqUUixTY0HkKVp/Gb5PF/w8UhbrhpJoM4zTpEZxM55wJmB6kv9xaIIHaDf1ZmbL3/
MPTjRsyo1TKNr71CIApbJPDZMfk8rUjgCt8Ax+indvjlAYwnvhDbRY/e7CTEwVEnXFlIqPXv4+qF
ZcHyeeC6MleeR43q/mSC+YDb49vOHRc+1/yi8vqMIK3DDUJBtUKCQ2M0W9pb5nvuKXCfFwQNT019
nZgoumKZFQbHeBrp3Yn7d86r25PuG2GaqzdIHcZtauyVx/tlxP26tmVIvA/QItB9kGIa8vawHEBn
3aXclPu0SZ+GlvfqzY3EjcnxE/iK4ntZ+CtLSBWso4WdrAyybwT/03iIaQwWUePovs21XcvXh7h3
MnJbjJEKyJRxmIeTS9loKC+u1mqem8pE4wWl15/zuu5V3Rd+RSv1TN24KNn/CpGM5D1KqsHgF8Nf
LX8xcr+rB9zligGqXKvrJKJ0ci3zmlR9FQnHfUZs1cPof/Ixa59pYkBQobEg+tuGI1kSwer65reT
ydIzyLJHJS3CkAm6wNeJ3EzWRYdg0HnHzsRShryrgK1yCmo2OT93sWovkjM6aT+1vyCSILd0cw32
8vdRjXupBdh9HRwsxafb5m/8I63f+/OHaJOYYFMSmSjo9XL5FEGCQJ9D7ZVMIX8duCeQJr8UC6TI
RpikiXclZoMaonoC3KrQPBoJ43peltIXKrudp+XW0UCIoyBNrfD8hpIyvUGtEyl++DZsWJfmI6QO
oQIFeT5xDY2kXGBorcUJg7MiDv6LLmy/qObOYiZZkiFwwjzYQyegwb3C0+u9F36Rv0HOWd3SQ3Em
YB35CiZxleTDXji5Pn0tUR9y0pUeeBLQqS5tsCU7FTfvF2aFWZ3SgCf1w/vXHllZ7A/O3AdBW6Cg
5nrKA6pEUE4L+nHqFxq/GhbPlI6ytRSxDpBXm8DzjnvM0k0ndKFsq5d7tphexBtTz6IR6/5hrOpX
6NS7+qN5rgIRZPpYUF0WrkJLLbFlpgztLoaYLgrpFFy1n7VZE0wcN9cuwxt93tGo69hWd4hbZYJl
GNUBs5oi2hGVVld8V5Yc3mYBk+l2WKPmVgjxnJfPaE2eZZChUYr5UxzG0mvfPRBZC9i7eyNAH86V
qtku+tGj8AYPgXzLevHkglhIwyF+JyRn/4K9hh6OD0r/WmgDg/tLpbTrycKTAK3fChdlIbWDLVpt
SppYLNB4cFSu39h/IlMXoseWQsQtRVLosXvdaJzyTlR3Dau9wIbN8/BRoO4N0Rw5iARDiQKqJQ3D
ZHqOeEa+dKwsddpIjImHJb0WAC0LFy4AFCwvbmvqcDlZIrnylAx1u4UiUFWiuHXzNjYUI44tM/nS
oyQMz0ChSnInMP5nsJ21sHvtTi/kfjPR5VR2h/eOiLLfxTMPqwiZgbSSuml7iGrpXovBwdIeMgMS
XEQ/T/ZK2ofdC7XIu8tSQi2gDK0pP/inc442CbT1DtrIrViPsquChoGkjqnancOWXogB7IMHDj/2
VoAIe3o/dCboUC+UWChVtZaYGnvrExqvBuaVRAfjILc1lkkltBN15HnY4PQFIQ20lIfdgPkI6czJ
lEryX13MUsXs+s5doQ3OpFp4+MDJFvdiUktFaelKGohEgnNmrcTDPyhVsLnWZZHu+EEMvqgJkTVS
vii//nsVcoNf5twjasktMh/KB/WQmcUK2FbtcftV5vQ21fW7cI87k6aSA9J5XbuFATGlXBEPoH/u
T/MY0IwX5UJ+3lH39NhvET4gnM0Udy4ZJ/2e1X2I+wNWdF9LAjMijtK7ONsXM+mCKhPXv69ZCx09
PCfNiVJ8BsenxpWHMQMNdzLOqokWP2BN7Tt1bjD2AdMACZlhPwRgP4xmygFpzuP+dR14gJgxT04+
kfTQ7i5Mj7aLw+Jy13enFdktXQSP5xDjapnNPOfD5iK/4sz/p/jlHx0AiDLGNZLq58t3O3CpVgxd
euLYQrT15WHKNB36iKtQoeiTEEKw34Zmr3T0bQ/e9MUGVspFCuaZFwC0nYh2MG0xTa7hD8Ixqxac
JGfXjNpSoOWurYjzSzhj9+Ed/CRlqZW1fzVXn2Y7nluPFl0azDYgITEu4K9JaAKqL7eSGCa5sLjY
6l3o+D7H++QWqmwaHqH7PhOphDuPhkYggz6CpGUWBrZ1pw0d/FzlP40LdbW+16qoZ++0dLDHmVaJ
OtYQW1alFPUNC1paBUY0+R+s8fVl02Mk1rKvYOKUlo14ZuD6D2jLlbTP/vxqYQcRq5vBXS4wtz9z
iFpQonmmPSF6YKRT69uft00wSZ99lKd0LeiCkZaZZSgSBRTC3lwr9KshmFf5YA2RPMExy3YOKJwZ
EZc09hkyNS0rBNpglz9MGyfiTVtGMoso8iEGGHzU01RceduWUlSWU3UySITUzV5el+icxvd/tthw
blecmpCJJ0Ivt2wvmNDFdMOLKz5Wm98MeZWx8ERNnV20b3tjjDDp8gchetZ3aGJiD4svv6m/5RBN
iGXbOjp1DRyG5xPHNYrX823h6Aq0sYzQY53kJ8WKEp1LHLWyv+1wR4Jbmv4MiABM6CTHAqwbKfOB
rBxFeGHdbWzf05r+hDTsnOQW2ouSpsGvQnpfOSmS9NF0PTk9WHdlL7aZN/brortrHSu/uxsBeVvE
5kLhouQO/mr2u1PGGIcNymuwXKGZOd6ggE5OehOiH+ZgJ45ILHiT3FuJQGZd17HN4pvpiJUxNhS0
HGTaBJrNZs8EbIhB28kMnO+WQbLnY+1TPfCOu/QTKoA1Ea072Avk0zz9PNq4fnycKJV7cK2nlqsx
nDJW/mZKWmapkqo/upSd2SHNzZGpbDdoOwY1wY0dpPuGN7SBuSG8Tza6Vmi8G0XA1EfabWLbdpGT
jJsKq+PyN4IOcLPy4Ogw+uJZSWOqfjXe1KOub0ygcgmZn+F/oFeCWcVFBft5QjGrhtcOtQq72+0E
hwMmWCm1URtWbL/fs+8omstejd1uA5WQ/2+ovk/wX/BKitwHWpLFjaTbkOIBFjHgIefIYQ3LI0y9
N9gcYO6QpnLyfsRGTKXEAmFUx9R/d1iUmNFCon+ib7q0Megurdzq6dHIqTQ+0PK+Anpx4oZ/TgBq
LizKnOfDFkWS0GUMchhjTIrRlEZI+6Kw3FbUneVgopEg3EjadCWGTETMZslIkQVaXQSKf/+CTBg8
TEZMnhqHzNmtGGKW+ytKlQqUkJdB+TVi9FQpoT8/7DI6no0gLDCI+NTHxu22HVm8wnTyivQA6i20
YIwE+kX4yQu4CUHf+z1GlvEH9yFpB+qoiE+F1MSg0bSyotP2Crf16zt/rajpytTNkf2Axt5G0SEm
bMAksXwl+vW2+Cwr2lsYf5SXC578vap7gaOHJ2966zGI5YSCA9Fxe45NCSqI0SVNjA0QCMIJIaAI
H3XRCmDv0hPzqmIPBokFtu1wPcWFE21pSNBZC+eh9IrTC8cgeuW7eOkSVeMdBdaFuYY1C29X3JdS
cyHtPbUOxEPVX28COkK3PlLOgP5F0y3FvM6jFDjAtHPWEZwjYNuDc4sE1MYoEygdC98MmhkWO69G
Mt/seL7NO/lvlytKySO4WMg9b6oWxlEQ1UzMau+H8+GUoA+kmNmwDALl8Mmvt25GTNuIq5y0DtF5
nCkpOXAA+8RzI2V4f+1s7kA6y5WZ0WqKRtQL5yTf2FYjM13kYLSXaUcruCX4KZq+md0BLx5Aou7S
RbeGwkdUt7612sipBw5dqgHdozYx9oLo1Ww91Ch9gW7DYqZtOXVEyDoXKWQnFJ85VLkSHRaG5c5O
2gW6NmNW0G//26Ea2uctABzdJ3EfOGB1w5gosVucCVjGlnchfFnAiUdDOkCgdvil3bl6DoSgjeBo
EZ8/1a/S1tj9Z9zjZ5hRR0z2uCTGA260uto8Nia9FbSUqrVmDDsFAH+HtZKY5EY1sqWkWrKPEXuN
YzmrD2PPwN5mVzI10yxXJEWcc/scCP28rbtosPPaLBZnAwR2Z3KqYY+ijujfwT9CRG94hczJAh+9
0u1wcjcEO7oDDCLCURFKCYNXHLt/KipCFy/Ce2z2t2vcARJ/qVRRi4I12iSdckcH4ECLJ102pmtw
ukKY+hgz5QG3sa1gqeqCEFDuQ77h5VeK7WE0x388ShRW2y3VXVqln4fF5hu3KCBN+lENFEY6ClUd
GnYnp9jZWbrHZIbwW4pCYzcgNyqeZt9Qs02W9D75kNbhgohnx//0UTkZm3O2EAuofpPPTxhcDYVj
6BDGJXQ0EA1EIN9JITB0DLPYsWqkZa0XyqEjxA/TYJrzHf0I8tF3nsoXgAAz2KMZvYS69ofWkJmi
L1hg9+N57c/Qh1ExpJLHBJemdmtSvuubd+6KBSrj3khmco5SGsBKM8opOjy5hCzwqKFvFkzD81Rg
40oQ5KGPhShac98vzDqHw6DmgLKd09mOv2O9LFyJjdmqCFAycLE8YQLIBvUAVujiKK/3ZMa/bpAf
fYKdb9qL6eaM3wF8TOluyzY/t9t6rvzI1dlbGVcTS39BevlXDA1sxsh2ki5ht2qvUV2zwtMztXdO
aaMRkTWCwhuP6wgCDkq6GalfJbCLlLkzynnHa6s0pPun7gbXyii4h6f+2jAB1zJpCP3pEXtDQYQe
51N54a4zP2CJiDxkH2o/qCVpNXbxNuTKXgG1od5SBrLW7D/fKVL3dgFSIViDJiQdiiyroWjuw95+
fuLUJmLKzmHBwQ0DTggxzSQv6pva330yRxSexHPfZN+YeTx8GWTtSvNnsakBuIbR5t4qbh0W1Pgj
9y7+H0t7ps2v54yKF7BWgt3E8XCPvLkmI3+B8m3oXlHRoEPuoimXOyWt6J2hPScj2SDYLz1I6jVi
qOkInWYxRrEdazD4AXDBkNxIhMr9YOQ6TbVSw9vuPYJq/1L83+wl2v3mDi0MqUO8OFbG0t+8igN4
I+HeVoChVxUHPh39Zs71rBrPNykaYyQx+rlb09vI5DnymcTP+EN0EbZGFHnmrCa9z1OJNJZjOaRK
tHt8FgaEnKi199j1oeVPf3rIeRhQTfJEkK9LbcdQo45fDIwkyntoszfazYWV+lK1geAPbRgGKl93
Rzzvb1fLNKBehqz5y4A6jHaiLVXu//4Bcfs4Vi2HJmmVsOpR31OYXYtP763bN3ccavKaVbmjHxJN
RTQs86lqZKoIANKcBpNF+yMBSoWt19LhAoEQRYiHJycHytrQKHWfjmlEOOpv1YtDOLzaht+rIiqX
bj6ILqGtegNkB8C6dPiuMz3uQBDl6s7PytUg78V9Gn7h4ntr4fvR7QfhfgUEYEroXhy/8k0UsodT
JoIT5Cvjy784zQ2f3+b5UK+xo2vYBVHu1RaTDfZcQx00ds1mrzUABZ7/K9A/xJZxzB3k3Xg8wR2s
DNZl4BSnvik4uxgC9QkbF3UhstItFd2qBFdCCD2cQ3Y/N3wChF+E8cTheiu7vl2+sKivfLAnKsn5
kcPcO5eaBATlMKdm1ILOe2rcGmwBxGSMHxU9YHiLeMb7XsZuOF2mvd3AfsljHwI0J6XJaPo25/3L
Sgy3vKJiEvh1ggL1Z1twPaF9wtHBo3jGgHa5SCQrblW+wvli89YTuW3T0CUxWeodgMdptPXrwN4e
+gTQ9dFrHr1g39B/tt8Wu0uW4cjK2H0DZgyOakf1NkrI+3iQcP1PBIslwnFQJbFjNA6P1JavEC8f
mF+C/vwcloSwjpnpJBln3A+/wfXLiEPWx/lmh19WawHlpd7/2P01WvArRMDtd4HPLuhGt+V4vqXA
TQ1R6oRs9IDR28Bsv3iDAYWQQgFw3PbuNftvKFjrY7CL69Hu9dCZjmkUMmR/FRvD1psaWFdif56w
rePEIDzrkh8O+nVVzbb6poHh4SPHGGXPxl95mp7fCow6uAvC4nc66JgPwKPhkl2g73AZlX5S57Pz
kjqKtP/v6SlTfgF7zdu0AHucHNRVRX52Qk11NCO3kAmp+5Gkip8KHPRHON4ccT+uBMticNw1I2Kn
LrCnqvKSeJdR3yFu2Aym5AN/Sv7fxuYGBwhpAswUPZxCa9Q+dWSd82ysdpX88hTRfjV5oAeZa+e8
7eb+IZM2ivPo5x74Lhs3ZlNSxU4lsjGKb54CGjCYO/N+800wXDkM3FSMhLLeEeAeTyShUo7fIqfI
QtvY737zwtvZ1D/S/U6p9UVUVaHinH/olrFZEnmg0kfMeLOLqAiSVlQbDKmir6Q9IxzYBM3tL6wV
gRdNgH86VQTLH4eTslM2ciXTacu1dssHmoBiA5/dVKiyUozEWR01j+dyHivTpFrq8u0i03wRI8wX
44LzjM0zSBtPWv+a+l955Fja5Bp+YjVQ8rz92+l6Ksh2dqDItSgq9xHQbkFxxVq1bDHhqAnBvMe7
CiwxdWxq2coLuy2nsu4FQHuXte8Dyes9C1tJZlvS3xKPN5dFyRuDe5+AvA6V6y/WkMsg6Np6nMKz
y5wQLJDzAKJ6vX4flPWvzuK9wF4HCaSbOcUrlJ45vbPIeuvyPC25oW5HcIcJ3V6xCLHzWGgEF9qI
iJV3SNzuROG7vaMmuiu0SBPmUP+AJevZibJcy1vkm6OHl69FGu1og1DzfxvKRrexO3+oepFOtrX/
gtO8CLfQl/SHpjnF5pu15/ma3GrNmSbSZS/qWaAN7nH/zT8piQHyoLUeOTVBcH4LSQQb6gxTMbgO
uQmZdPxrKVaLk/qQRVIDQoEphYQaFV0bYODA/dpS0RG1IPBRNOwIPacSAmQlkGalfpoNmirDZQg5
R+x+BaJFhDUSwEzR0cS2zsjwt/F+Muj+IY0GF55ppJ1DElFIMl8m4NIl3Jeuz9peXrwagvah1qqe
DqPaMnl5TR/7phoX3XKtvFfq1Mh5rtObowRW10q+QZ6k3j9Vo56wYP9H1eze5OioPhgPOJh2ixQZ
9AhJR6WmfnQr4Lp7K0avuuqXA6eVoG6ydTlilj9IG0CsYPwRtwar0eJk00yh561yMhXECNpJnLks
TLDjazuPdw+nOtvbcqCkX4O2xGbp2aRbLxCfk5I2T2mf08AP9SEpvhdnykH4IJjz5ihXzMkt8CD6
pi+VVsS9/az5wkZSS2UIj5TtWZxf5iJXau3iXh/3UVqFCjd9iEWc7eozucU/3xf8ZJGxQruIu0A7
iH6ibFF+jN/kUowvZU9wq9AmE+RoXWl+VZsO9rOhLmDA6nmLPa4vPt2L5Srszsf5lbnQ+w6rmHtX
n1ZQL6knUe+DWzz4HXTXkCHEkVMoWbCoD34ImxRrwyRvnOZ7jxHR1fWiMIkCriYt0eBw0QHtPUIM
11UfWbQR7z7sZPCmCyBQ3MqgvOEI0QbrLYbJpgKfX+N+/ziC7+Z0h/7YEPJbwcIyiMp3LUdW4pj3
PewkBCJ0QY1bIjuiixmM6meu24Que2v/mmwxIIjPgzkmaNg2BuhaqUdac+MVqJg/Ov5/5+0c+7SW
0AhNKLv0FT564SYt0KhkHKv4PSExfgTrt83J/QapKU7Q8DGWTJJgqZelXmW4S8qmRHKhyEg7iV6j
+huGFZZjhJiCyzy2upYUdVXCYzXembXrg9cRUe3MJfsp1sLdCXZddHqepAdPDespDMql07CsIsL/
jGkuCFxuoUPa/Y8zwDsQc7NcVZNoetWApKxe6C0Yuuafq12hn07m+WPbOyLqCwp3ZxhqN44DJLkW
epkpn7FT8/ZEyQ4+tqLlo7nJCG8N2OaMsAr5pK+83WFB8vgP8D8Bi2gG+3mZLWFpXPeo4O4hlw7z
ilpH03pDKXfh24wsDIV84OJYKhDABm+hZem81Wa0LiqX3YNi58wELuJATegiYqD4yKEs231M9ZCe
/LW07WlVBbiFkx2oqxDm0zvWAvvAl0YS03FFijK5cPekvRGNI2UyHt3s0JhU6V2vG4tALlRafFFN
Xq8nhGdq0g6MgVo8GbmFsSx5Vlwj+leQFek5swIb1WYfNKcSAJzAsPZd41+1KDVt81Ha+MEzzQp9
k6vxhHwo278VcGtbR9d+CWVzuqRrBV43wRKdjfh8w01L3K20sLUGY8wxiPSvkW9t2jtYKGaAZnFE
rwTSD2IK0XPmB3GW/HVe3sgP6ZRptRPyC4W//H1jT2NiMsF3Kt0+bsXfVCoV4CjOB8ppWky3n+iy
Ox3KXxXeG+3lrBEiw3X/Eg7QpwhrncKapebi2VYIQgF9JfSW3Mjmi855O0sZ8jSs2b830t/xear+
aYyb8hbZD/rB0OcdIEDXmt6lWezbo/VTKSJvxWL9qvOjUHiHY/B0eBt3UMJkSyiyiUN+1Zr+qWXR
a3Vft0vz2xcQQvnfy3+Wn5zL2peJnx3kjfxLkverBJn7GnDWkak4qAChdPlrHW8O82oPmWXwrbiM
ab2bC3FD6wTjcFo6ZedteF6micCZjuWMherRWfOC0K3olNHzoDinE1tSRuRFIxxB192xm5rdmCIq
1oHpDSqlndpWWd55RKNP6B9dCxBclGnte9YV8+M5Mz0rrjbZ7riJU2/sJ3HEPkvJM17FNbaycxXm
uUPAfq2wAqKGAZc/UceE88u1IPStelLVBrw525X8msUtSRyjxVXGRyR/QxBuDFjNz0vJJnCvQppe
T5DY0wQq8AN8Oyp/of3P6mEw/kjadEEuPE2Re71oyISNr9prNB2iBHUIrbup/LbhoAU7SWSNa8eS
FUP1hqMQmlCfVEg/d+naOlmB6g5rqPSBD5hWDT0eqsjbddS7gEGwL6wEtR8SAoIrOPpXuqKJBaFd
DTniUAlpIt7haRk5o9LlWTSx59jg33SVW8EzkOIqm8W3G7DFmVfGxCA2a2q5ECTR7WrHmqESYaIL
uylmZKlsgYZNFmpJUwz5mt6sgKIF+O3eKNT5lgNoqXq9qSiGBaUqA2s/0jopAalyj8iULdF131RB
0ZCkmXwgv4UBm+qCM4RhMRwjqeLuZ7N5O4SrEw+XqKc6HrxxlptkgFNtOOP0O95oa33cUfB78OEu
AKZUbI+XILjafEjIvcaxsbYJLsP3wiH2+uHr7W6ea2Vi0BbEKboCd7kCPU/arABDRF1c7HeaJeFn
FtdlZDgYdufMKVICqfwe8MAPlnkEzI0VAFMojFlPlWTp+/9J+ovz/G+x8AfS+Rn2JdmKjBtuwlDM
8QN7aIq7hFDb9MK8xm/TDJsxQ/HeSGDHpwmoH3+mYQcU08eBQWgP0/X6WcncqcZ1Upyl9ilG+uzB
c2QrYUEkL5mBPX2jhkwn2Rl7ZVMNvKAj+gm532YzzTRVNM10cEIYmaQYDoAE6asNQbvMlqD6i2PD
PNeWAmmNgQ1L60VVDBENYUA2LtIj/LoWGkjNrTDsZ53sDWqUyi4CIXwi/ImBip4JoZ+eC+t/cOP7
TYOUsaJdcS2GBEKTqx5TJC1bYAb5J1p9LlxMqzj8hHhSid/KW23TwjyqKzm4Ub9xKA7+vPEGpC7R
XJ54F6vrICHPXxLIeCCdziTFJJYIfetX3mImD5ZLlOTHn//JMeFW+OmLc6pUsy/0mBmbedrob1PI
XKnWqmmGUwxnYMwackYQ/B4Nnv/Lf7q/7amFoFgRU5e1MOYEm4CVLxh3ngjlXkNA6VEUIcG7Sh/R
LERks1MEXQaZiafXs9ztb01YCaDGA2y1wAmI9/puLI2szIxdfUVQIvyccDuQ90oNkYYB2M3ECyGm
WJhC/fbnG9fNSdOvFEWcJ1UxjYOYTMKvtqiUlMv73IZ9s/LlHY2OYxlwodnhO8WS7gNO0+GT2IpY
2Yinpu71/tGlsoCtUYLosiPkDKaefnXYqRuMxaw85emMR1dJNTntXSpGU+Rck3gKBg2gVTbXyv92
ajO6vhLoi4FJwbrfMIypM6HEgk8GKAOsd4WtC5sQWdBIzbXnIhspmAgI3RuP3ek/N0EbM0GJpGgE
y4ToeJJznTF2uG2grrPLQ07PQT0fwUAdD4LLAE2OiY63zf58X4TaKzHYyBgGag4hTeYJh+Egcjyp
MCUGryjoSjp58NZOvIPoHSCQDrEO1N5KMG4O7gYdQikLsDCvwqfvbiyX5SwDmEWfItWrRzrQe04B
nkh1FA+1tU/wxzvO1SygvStrZ7MO4apmdzBqdqcTb/0I62KQrHFANPt7XWs/GcU/mHfgipmI8bPV
6QhWVu9HuaqjUcLZzKLtwqugmhtDI2diwWIKONIGllY05oAvF8uv3IvuqK2UUQB8nWkRVbjCKYMA
TK2SBE2w/tb9UUM5eDMlICREt/CYHUIWqIwq/pmTMcUGouR5ehFtFepHLYRAo5iyOqfPscGhSQmt
Ep2oVdPhBWqwW71Qt4cqzxJqQ68v2m29DLBGhMD2G4JajJAmPTWnptJHOSJzuWvhWi1j+tzfalWp
IbMcbiFRTQbVNVJhJjZEM+O8KklfeuUVtY2ZbTHzuXi1BXCqvoNv7w9xw96WdEhKYzrrZ3bZezQp
3X/dw4eWEnWIapzHwvC2KaP2LZOy5Wk+kO8lXBJC4pesWj6foB5yJ8i6SPlc3z4bdRqi0OeohD7Q
hK2ZXwaQiCI+MDl+7p5Sfrubc1O3uoCl0XRUF5HmRSjXKUtfSdIwEep7ljcTixkvULPBGZtZSTDT
h5wd2ub+zw2+jfL48zALCmpOIVMsPq6sylkDZ5o37DhACcyt048bR1Iozm8Aoyo1VIkx/y4RL/9q
3GvgZMa3BE/DA3EjN3iA+JIJIVLK42I1lE17LwwT2G9Sf1WSiX4W/2pVUntiTgRvLPPOMNkQL8Ou
bNlgI/QqSLysLgDyqfvt+JaGng+tvYK+hJtVAHJNEKFZ7bsZZOA42BuWI7VGzWBwG30YKy5chY3k
m1PysQaFnGvXZQlxtxnw84lAVW0vtORyeykL5wsug6b7NvSZUTP+/D0wa0gyNxaq5mEm3ShkWIYp
ddRAAYl7HhS7Havdxt8PUPB7LB5SZqCDu2NPxNOP39crBKNq6pu0Gtv8nlgpVf0usZeqz+OY2rZZ
ALgOsi0n83teq/NEpW5VirgDWKww6MM37mKIedspz2lU5xyIb1ellOhaPRdyGN75FDgZ2MlVEnZz
907kC+x9lNvPEfF6u4xav7CMCMd9lmQotAWNHQzGPglHEjJCpiqM1o8wQYBhlJztim4SVKoDWM0A
GraRC5aWbIL9kX/ddd9cyxl1TyPc1jOWwb0fiWoc8UUdsKO7xAJdroLGZeADFi/NHZbaDSN2Ob+I
bZc3QA9300qs4AGsXXEODw7Vo9U1F0n4IF2mnoOEihviRQ3KxXJ99Iwu/oSDGi3YAI6m3cEcAOcG
cbsaxRk/YpyplggjeNe5oE6wtRmB3G8D/YFx1nqtoUwxlQY+xXvTk7PHGBwPY6CboYfmCHRqDLqV
qVz2HFxdL51Krbnri4L5YgvuVM+DVvOnpQ3XGr8rBNcMUxf4ZgDVpQfOgFUxD5dk0ibUW9v3S/rl
rGze76KQ5LZs0M+AYc0pW99abF5YhjcLI90DSc+g95JdkY3pVELUePHrDMGpMus6k0Jk4pzmfXij
IvSqhAedCZhwO9pFKPprc/BjYHqWzjiDQe4wHJmbn7J2gT0XTdtS3zrdthAvJLnylWeHgVviPTno
z4TDr671kDdG9aQNl6CQmk2VkWj2tWIZ+k05/LHOPWlhN7eC0ewj182NrVXM/S7fkme3h0f7hpdi
I8g9MSf/8Ro7GEtr0D8m78iReQlmLcNGuNFwWdEFXclf8UhMoHenKbN58/VcjflxBlXCa/riV/Kt
bxco5IZ5i27SxW23g2hZrKZgfoOB/Zy/cUVX0iohllY7UQ56+GAbfTc0EMSpAeiQDciyJTCaM9oc
equjTjmREvP2SvzXHB8hiMl/2c4kv2rGOZXmQgbeSI5borgZDtrelN4TYYWldFdQj6chWUX9lqB0
gMTPgBOsdyA5lJ99yosRe/NqdQvPOdynhMoq+BkYhlSaeyA9UGMb+43O7s9DC6HTklgQrZCEEih/
OuKwEa1YTrlcYqKNu5rTnTgzCVWVIxdw0E22C5GM1If1o2x6y+7G9E2p2k9coqzO9lFI6V3EiQqY
lWHXF4Uf228iGtrQTkppO0n/qgp/ZiOj5qhZAz+FA6xCaFD8PIN8/ekhU5CAn+56xD6kUbSx0cJm
WQ0hNUkxjVCNRNlE8OHnKt1wTKk/2v3+SoKOV2j2TeqPdiVNLIYvHXk4UwFJuL/JnnMHohiBBBnf
XY8z9PQ89seVti55ouea23//JUyllRifchVADtJMNhSeq53a3c9lKZws/I82MQddU+ZrxPrhZY3J
3E8tV2BqRs6/dSSS+VwyYMeEcRnpzinD8tz/bAH/7BqlmbTlJ79JUsItimUpzuHj+TzvEB2AlzEw
PpSba7SkgyBrXHxmz/ZZ2GmSpQISdLB9acEmbbOlwHocVZWYRpS2vcYto4K6zsL3M/8uo9Qcmsbt
pFGrg4MaMR6JL+c//7EtLnb9XjMtoFgKilbC2G0kCjlwFuks53sjjmPJyb1lx1OZlyAOwZ0lPkCv
lz+98DeJ90vLKM2ZxiaLpLUR6ZGelIeENU+4iJ4lvrmHjfv1kGoDjS5CAV17uKDwD6K230VA8LSd
MBoAbbrkIkl0FnKCHgrmjslhllYKEig00K20qP97fGyHbwHl67FKGEd3Ny6ur0YT49AfOYhGVpJi
F/HEnu8YYgsqCiFcaBdB7KxzD7VD4DY4F/bFpmCUKVY/Qoevbc3rnOe4YsmOecDG/EsY6z/ISqGH
adSwH8I4qLjra64TgjZbcz9qfk1yPkCvF/0OKRmuPf7s1/d1VGfG3GHnL/ow2dJFG8g3LD8M7rif
MqawB89hRpxAyDF+WQdJtMK+wxh01r1hEXVWjY3DJ2Grmc/fY1Humra4qBctgTYfR1XcUrCG+//d
AkM+CedE0EB/Bxm8JRftkdM9OaY1Mmc0jEZzQpSw+gbcT3ebggbAFacFRECaCUTi9Zxo+v3q+lle
5H37zgG9vXad33WrKS9ROLL+rhDn7D+QMFycNJUG2y7kFkoPEq+95hPxDCObbIL9HpXaPuPKAkKB
rj89xQ/gvtj+YMe3fJBKQa3iTPxGFdQVbGFLvbZCATjJDFVSN0fURBCbeIe5tsvjcV5Hwq7CeWix
PW+4dktlUvN9Cgcv1JsNsoJ6QYJQXVOJ615/nTZRpH5UFIPWcHSUalSKUCg/MW8LJbeccRm5zQlk
WCm99UeAJ8KH+4HWdmVfDLPvlBgulZR0Lcl1ERjRUuuucQOkTY1LeStx/ZH4XDtK6tXSqGpXYCYJ
6X32BFdC2A1msj2vbQLoqQjVM1B87DqbJbnbHXaCROCkAX95ftd7SuCHlyb1FNF06R5t8QNcU4XC
Pu/mckbANOF8o4v6bFGHlPjpSA+qJ0d1G6tXEJj5xrnTd9IVAWPfWF0y29oqjO5gXRvAc3JWTyhA
Q1WKlf2T7bbSBERYbFBH4rW+DNWiDyv2/Za/v7Yk+vJ4n0dOLSREftE9Gn1aqowSadigAhUyNDPB
/9Z8+NKzBfxAZF4rPeb+hywyOz0BqhLSA6MeG6QgASlfhspI9gkV7pmXFuRP/PsRxx63yVYGdE12
uLadpZ7k881tSptLyXdwN7cQPNeF/XLlLgSot6V4fhgDVgtHGculifCxd/mPDr1gxINvA4kNGJUo
B6exSlrgdLYYE/7VNx+r7Ax+I0G1HvEp5N0JdUJpTfRJI6JxChM+hK3xzbVdLiplI1KQr03RhcqY
lZgeofphCVZXdjDwW5cZ7cbYFWjanW7fhphQYjQSK7L2aMjNMR11wRyPPSf00WO0QT5W50Xmcw9G
7ho4G6z+I/yDVU0wGUMbAqsCNVTxssFlU0AL7z5DcRvpyQtYMKL8OvfYqw8Mns88JhxfTeJ+UONO
9csNqnm3ZEY/g3ufdRby5ibMDxAZbQgEVEftQzj6wqh2GMWPD7wmvk2HNKittMy4Xjfnp3MvJQLi
Dt7sedNPupx4uNenY351ij870KVPY7oxsEgXu7/oHEFze5t4l7s4SXrABtsMw9MV7iUXJ55JweWy
YXx3IasAwpSejnspJ4qqn6n0KfAuxnxrn/fvu1OVnkS6hYsrMniv1YEyOt3Lu3ikLFrTKnX8Sj0N
jrGCEnJI9Ws0/Xtt+5e2bTk/Mhs090yHGDg0GWyeT07AZVI7CmD3clYEl49QbntXQ68VSRATBcCB
t+yWTC9eiBMMSYfqvBzHQCjZo8L3N38jgU9O3VSj5t7d9Y3n6kGOqghsVowfg2omjKJgXTefkJK1
0N6EEMvOz99QuFDgrobTI9rx7nVkvpup1zrotBRFo+mI5OyCP2Luv7ob2q1W+7L64QfHLWBr93fV
oekhXIw/cpvbOwo0OHwKGCA0pJO2+SiTncmTcOILYXwemjqp3wNUtRwkOqjXlEg22jnE7x8EHHHG
IIMRnzRTMRLYuywgKo0c9om0U+X0vTUw8ZP2V5Ziey0SvSLvDs9u89cZoxRdZWJId3kXGFmXk77K
kQhKSphXXwEu8uxlhOZTOhiByCFF/TSHpBAyGAIKTQ+TaqmVfO9cDbOufoF9KYc8dvEz9yNKG9FM
NNr9D38ONtbPFiRdiHxQ40e0S7zYEHlByVKGBV2LtwULijU7rWuyQIsQfGkk3dv6IvHyciZrhAJF
13bpu+iOljfCfhvB3xHiz2Q0J2ivgRjvVhD/YuoQltMrvLBIR/TLPUvTBuvOtkdFWqB77nzM6t5R
qpe8vrR7ZhGFyCgelxY+N3oFHMwAGXbRsOMEKkKF+4acmwf3b27ul7lx1jlRwpPhMqrkQXicytUL
sXponDgCDU9RdkgkAQhC3wY/waxrNHlVpJVkvraSkCF4s0HOfS94Fa+hm4fDzZ75afDbqkFvHlS6
aMBYRLeyM500M3F7viG/iyK3Ib4Rzn4utFsdWLQ4vSTmDMJ5SCc8C2btkA8oCqjfb1YavRQ5WUom
e6AmzprcgMDgBVaqq3j8kmZ3lGOlkbmlR+qJCHhUDGhAnlSbkat211a3beFKArLMQ2xTAP+aQXyp
o21MsiWTmh2C1CkiZkq5S8VIUbyrz9/d4dCmCK7nmVRGOV7KtLodTpU9X8Zq2NUmP8IRKh4KR3gh
qgCV5C+Rsk71QWuhxSSwuRaexiYxOQev3zWu9NAX4G1T9uPIycbEhf2jGI+xcoG7wWBJH4zaF5sp
vRNWb8MXchc6yeP0iR+6OllpAou93Lr6K8wmb8A2WEQC12XeIQ5msCBmQ/7H6iXZv1EU4kHeze1M
W/RrKXYVkhmc5cfR2/7tde3+hG+kViMg0VLkq4LY4LlMWimb661G/ter8/pWevAqu1Mzm2J8FLci
YkNdA8iK5d5o9Mz4zPLJ8RZjK4ZSqjDx7tKFStKiGWcVWqyoSlqkcsKq/9+/yZQ3jb+gVNWMUB7q
ooUim1jV1MYwmjcf5M9ipsTtTtNcXA5vLx516IczI841lawx4X5ZvLrKwiQFoZ7xAa7yabILxaLt
eOXtmMlmbuAeSh3z0I6BQ6Q0FoQNbv3FXROqS37cLKjFZV3+BAn+hiAQynqeygC6cU9+wOBQGKj8
fpVUwQqH1U+4WbiiVsr4q+VIygu0FciMBrigvJ/vzKXej691EPxhavMwazABTCKNun1Nz9l+ueU5
yOD7bGuZKd2GfbLvD2fqqvmsfeeJahrSrUt7xarwjYayA3zWcppn8xlV+ybA2Mb1pcUIHXdk4ZX4
0r50AGQU4+jzr+9kC2ZaVcx1erYmK+l+N0AQFip5ndK+z/v4c7MY1UkkVUYzI5E3t3Of5pKI71zW
QxcUCDwXXPmzctU0WwCzAxvvX8bLsRfLMbt1W2xgB1Cm7b+eAegxIxspeX6wecm+zJM9S4Buq6Ok
ysuDvRKfpCY94OcI1IWALx1gcAYccTqM79sQOfo62CFJ1Gl/ZMRx7OuuTHpfheKKx77TAC5pNmjv
FeuRD1ksB7rfPhs9Y7cKtCKh5f9DhKvX34lrDOcGZ4m5mu1/3P9f4EtfKTzmZvTf1eSQxGKqqmTA
vJnvr9fX06KiXQuIXJKFTnm+k0X0t8Yrp67BLmIruwP8GPLj7RQJu8tc9bBL9cFsp5RQ5Q4P1ASk
3Hj0uLy3bNG6jcdKyTuAU80VS/nlDIyHekgUcrxuhmlELpHVUIUXCsShLiX4sz0JsKQUHbJ+l2DR
Mo6zJkbx9+rpJAO43uwxL6uEcK3K4N2vhAe9Ut6mQKOCJFIM3ZZXFc2D54ko5Ji7MXQIdzyWWtF+
6IrGeSrJvzhXaZjj7q/IWDdKi9LGikcYAA+9OWqMqCoclfF8pVHJNwjpWr246qJwggi6DDRAhbFD
c09R0sqhcNCZc6Q/+9mGQhJQZlW9qT4gKWVAP4EuOWx0k2TX4yuQ5WiMb0NyLwjwnjNp1pej4Tpu
QreS6MjUYHbIy/ldzbz03avUPx6EXT2cW1daUgVre/oQIXOSWqkNz674GwGQ5cWkRlIDN7//Mksa
TCGUwNdQOTtqKotV4VYyrdvfpA+awfefHwDy8EVj0jICxRTSYCsnN5Uq+H1Vu2p6j7WI3mQo9SL+
CT0qodEM/B6U6sG02Q8wnQIscpYbjj4XDgWb2HUtJf577aytEqjO6HBO5nr0f8nsrlIieuQwQKxn
vcKyD7kU3a/kKs30OTIFm7OQVU7M3QyyR/6ElaHcjAr+EOGtQrDyehxGqVHk9W0sX7WSWfpmOHNM
wnJRrFK5H0UjwbJEtbtdnHTsc1OAiiUG9ZO6Ul6dJT2ugLbvSFFwJCVjMacCosRh9xuJMcAUEM5E
jFjEPTsIFaB77npTeoYM4g67zDnU9Zx1UFWhQYNVskWNv2t5a3YTl9gtSYRpiK3DEznSLFv21MAz
lFdsBRSLdu6oSrj+meCTPwSicWswAEw3vPfIMRDyGNASR2h+1onI86l4tcglriIngEZYDPGc5Dcn
H2ezGs3B9Vo0oKsmy8A562VIXugAitCNtB0uwZ7jPo9LIpFT2K4EmN5k6xoaktS6FltI61rJRQgt
Y6r7kupq/1GycRmiflBfMuUbtkiVsRvlfdRDczzzB+R2jb0iU2XPzPiLc3XTDmQu7Ti63usiVuxd
JyP7FDpKkuNvhUQ1qg4q+qe1ynQ7OeIPypjjUR0BuYaYO+EuLyzLU3ULR2YFF94Ms8cF+11PYMnE
+LGHTGkJmvuaYWjhIzx/oHQ5vDNGaaE/v8EDUwUH2sFpZpxMbaUFyDGtf/CPpTZ59Cc0KB8C57Yo
FrPKp+hsOzYbnMbnQLiAncDkZxIiDQRrmpPhC+4tMs1Uv+S1sMa7+bPbp4dm56jRt1p/wGEGktul
nc1TopZ4w8ExkrxYB0OemCPY/WbQoJ1PWE4pz5zXDnYGkrFR3qfJ4gWXssu5qGs8lKIbIruq3+bS
9WbTaUncPVt15TVN2Re8zLygQ1hZayrCp7xbj1qfKQfX6zc/dSrSqRWPNza5C8TIus3jqm7aVc7V
J/WGCEFf1YXk+AfxWPMJZu8XDlsfAsjs9fFgg1Z3D73rPzUegf6yJYQTqV8xEvyX3cUwkuGuDXEM
TC9QXL5Rn5U20hTjpnrlsVC53RhPo2J9J1XKRA+PRkuGCp1XrNBfTY5t5prefuvDZihNBE8z18LD
H+HbgVpB+akl6nRRSxwTIEZa7bRF3h4GvAPscTVkP6KpaixyGTjVrUflF7ykIE2KscqXgAOubAqH
2ghua5jk8+SzXzy8Add9k/hIH1WNefmh18y99GhIEgn1bNuoOxl3MZVxSbh33yXBnWLmYEk0hnqW
RAGMeX2UTmOKpPE0XsoIL7hGsphnXhx+LjMmTK2BQaXwtS8I+crAKVwal7iTp5vq0n9dLG2GVCgg
7AXJGCwNPEeUrhgnsyPJ9n99RGWo98kW1snu7qCotrNeZJ+s5kMQjoFFBX5RDA7WaDKQo8cpNcvK
J3FX3bO7N1hNVw0+4sVPuKbAcO7LEwb9mJLHb+tWvZJe8+TzCeYqbIktRCioIKQfm1N/mg3TiwhF
6b79/lZItatczjklU0MNJn9Af1D1EMyAJSrgPSj/vQkq8F6wXHsZfoSM/EZk6cjM+FEvNGjbEPrb
rOqnEehi1TxzpVx6lClFWr9divHJw625Ol4dOuOuPfmXc0vqeUIDbuPMxeGhevek1nAusfsT5S2P
2sNctmu0Jts3UUP3ZSt3/E5khWJNl9errQjMSyUDLmag5enbac4Nlk04LjZ4dTiVtWlEUGCjF2+Q
sJru7ztHJweggPmKIjVHo9Ds6CYJtzRJum2iBMKKdXFNOD/WymHX07wsGGLxbggjvgh4NR1tfQQP
rQofzheLlIdWa7Rbjcya4fkYnuVe4EObMMqt//S8rGtVz3O7qXe8vJgnnmKUCUP861Wk8lFNfTka
R98phLKlj2VghRKky/R66z9VB+Omc2RiIGRvImSnn4GOnp+nQbHPLo9OvlvOGqLSEhC5vv9e4oWg
PbDaEEO0IveRoaBRt7a+M0pWmXaA1UBdU5cZuzoWA434625qzqC/aDvFc/GK0s8kzseTuoqAPoGG
tWTHbCO0pI2doJ/4Cm2PVNAopYC5r1xVDxptzHb9M4XMUrk3r/Ob1enooWczml9n9xaBAndHhcL7
OgPzkfUjVFlHt8nxmEE/ZNfLovXOX/e7tqMi0vYMqJ5sJ41ZQ0QvFWUa8mF2HsYKlKwxL+UxeKZp
ILrqDtlanTAUZgiqHr7BMBF4KWOsMLS8DqOpkKEcntccGJaLcBLljRBr7IPUMtj2ivyIoB4hYWcc
HxXUMz5R2c58tyRyNoAS4Pg4bB0ICemVt8+urLqQBc/tLCfpGlTAn/xBuzK+SbbtsJdfA9+B/Rxk
AlWG/8MX1KCs7I08aGotm0PldY6n33ZrTyzugcVwoS0B/HWbIL5UeGo18bsS0Dx+mghz4i2g76WM
jSeMtxKMnxUUK8tSc5KjMK150kaJf+EQpDKJ3FCCk1bGL77qTU6j8ymqpJoSlNFA+OiP832oUiT9
RZSNDcTdy4UNYwVEOJGnjCiqz68+6OBrvJK3Z8YZSzLzylZA7RHHm4BwBg6FC90i0XU+jio9viFb
gDtnbi1sE9G/0MTu7ePFGMywuAbWSlxG8WaMNWhXpiwYtLMaTfvp+mtioN+pSVRQgqrz24UQKcl0
IyXF+hyHjPD+oxaCUurrB+3SvojDWlYIo1f9oc4Eah9KtUGEMwZVMbjNCQvxt87IESx9EKIWVkJB
Hb/seNG33HqoAkpHKtCWvssJ1C7xjzDbH9Wiic3TFT2WAa2H4AJB+WKVbE96o7p5II8I+ZavA/H3
snFyyq8eN3aIND8SaKMGBP0IkNYzGn6t5EBCpYh1a8pI2KaZB8kmwKN6csVLckB6xaqDgmmcr5c1
FNwuUpvQ3jYdkb+ZYSCKcdTWZGv0jM32NYa+7OVjbvMNNZcVzgHDOaD/vjIJQnsUyzR6QOUCSeWn
mx/a8wV7lqa4IRIr6xKhTfkxQBh11tJppQCRyVGigPeFCXicf/Sm3IdyYA7s7Ky+GcWMDd09SELY
xxXJGOM4DKVwwaqxuZr14tn2wf8A5K/ka03VMqI4CoENDD4XwFJg1U4DrKip5hTOXiVY4hvhCoDi
fnhOV6+0+JVr2oR40On+RaSJRlDrKMTYBkhYzbtAs+SUGDAvqY6ajPg1ajhdvWzvnn1/PxwYQGjf
2t7DUJ0EeXckXYtnZNBLDm2qp9e4xuy9CfrSo6t3luMIoC4dMipyQeR6tsHE6OcnSTD34TDc/jAu
lloYQhjbk7DXitfVmW7y6aWKnRUqPNTrxnVL72Q0LLZWrfJkOFdDba+3izUyd9Ez82S6yiAUoeZ1
e3hVgYxn6V1YWGuTNLPtFai5T3zD417zx01/0jdRW4DYXJXxHEtemXHTGaHGgNnp0Jbl1147TR4z
JoXMZu9RDMlmLlU9EhsMU8J861j3r0nIEGoffrrB7Hryf6wVsnjR5dOjSjlpCen19ogPxxRXGXP+
WbPXW9fj9mjcbTAbHTn7m7MEBi+7rPOufIbd0PNO2t6JeG/P6wQrfUVlSS7B/V5I2B60AhHLEomk
67M/G+b/OKFE0IytHQpBIydr3iitYIsAqAz+BZYL8HFoDN/dYjreQFcStoKDOA7Db71BzcS+Q/FD
5SRfGb/sSazJE/AvEU4dyu0DAPA3lrhFhgIAUgoXyepA0Sut+fNHCbDp2X5QDlzyvCD3lU/AnpVa
NM7BGmkosVD2Zctc3fTjtdqsy+U4e9C/Haa5lan1nsJWvBn5lSMb6vW3LYZkhijV5b7Lk2Jqr/Uc
dtGMRYoueUsjYo0OS+Ab//kDii3b0ANUtkC2ixMWLxWHM6i7k3D1MegDmmOKDkHR+eQaofDbqQ/H
t/FvpsEWmOkWHf7l4HPN2xONAYUg60uxkCQbORH9svJABD6Cq0kroHr4mae7DqAZf+mqzhxkX3Qk
zLxInzaq1ZgQNTjdhd9Y2Mcr8rxCfBc1a//jX6cYbHv8VQYy8Dn69WQrYnAR284tFSPy85sE9/nP
4fVLTdgIEyUk5Y8ntLlfGc2QyMxYfOaktUCSfAbmSy3EGSvwjsHVumFYCMaa0lPGplXm8H/jT4Dj
ByRz1/mrzL9S2GglGERCaDO/t5NmONH+qbIgbGtXMDjBum7mZNy6t6zefY5RSSYTg95rc+XmOtGN
B72AhbYgpykfZB0Jly/jPpnlstMbY0jic2AapBLkPDwWMYK+FOi+XvEzPTy28Ub8vKxVTePP/O2k
JxxrILa8fYpkFEXuicTCwccGtLlO+qi6H9x+wl7vLiGTNrT7mB5JuexrZccOgExEK3EgSrRQTZVL
EF4ET3yFDidEmQpS7qooXCYNBHYXgV7mScusyP6ln2DE5gzJiRG2PbsBV6a+MU0Vpj8JU/aNxpMj
UTFcu9ey/jSP6eMPwD9/46/oDKIzGdZR/23vCDiDaA7RDUGncRVrxDPjErIJoEv4kg1dieNlW+hX
/fE/U8idb7zWZ4nvsQoPvLywwtjsmJwkqw4rAKiMc65GPmp1mGIxCLwMF0BzpHPcjg4qZmRY85j3
xLdUFrDuhTjEv5YThF7iml7DCIhJ2CxvS6Qkw1HEN9T+eNhhRl5A46KzQ5HP5nLKukZKxfczoEpN
5+l4xWOn0NLiyH7mJavyftoWC/JJO/VtH4/BBf+EwSnehfT1rFjtn2R6j7aXOgJCNNrq8kiWw0uX
4KqmvWRQS6rwGO9OoSOOK7Yr3wM+lJV42myMQSZj5JbEYUGj+zMWTZ9MB8FUPgElLc6moVB/t+jB
S6iLftKpdYX+1riZn4oVid0knuHPJISIwXJiXipLDe07ZTzhY94W2XFsO0Yd5SU6RdGssUFNF/Dm
lESrPYuDcBAlmDxA+8HwRyQIMl9SURvbdxUKCJHdPk0dAYlQNXzOMMN9nBrU+zyDgVDb/liXiuAv
obv63UQhYCWgf1EC7b4+nIFhkTDMwkvQdCrHCgpqViZ+dtmYxHezZrZVotnX8nISpY3xNK5L+QZE
CzAnzSbbo4CcqzETPOnfrRAsQtnozf6HQcA6pUggPJtyGuotnPmakUuMDLdLnMr20wgrBvososHd
K0f+kH64d6TayL7c81tLS6blHNHF57FvpfP1rPreYrR3F5zgSwjs9LRk6rfK8Ftd1c41iAzRq605
cVEpIn1mMDlkXkDNInADSpsKeF6DxIsCbq83fyLMEM9E6OuuiqATIrzm5oEigbrOhGiDjP5TFZMP
AQCT1GI8y2ijstqs0tfUsCBOufbnPqUVoT8kD77Hue+ESquk3G6EBP6I0deWDEHrHIZAErd58HAz
HZIOk+s1v4zjweGQFGLM2P/UbgLAwIfRx8ZzQYWcTo/3fyCyegWdgTgXyUhzx1ZqdYwJm1samBM9
F2s4dM4lm/Z6CPDwla3YJR+fXXQbpW+OHOeMzqC2zSVK0JyNBup+f93TvKilfZlwyzRaDzOI0QXX
Ds/9tqDrwmGbi0SJfKSMcBuR4uy5fShW0RbyzF+8W0tH6fpicrJFIiMyhHct0rpnTOlk9qNB7I5C
PekFdsGMsvds8rD9WMSl4uujJ9Vz5rdm2Jz/8CQjI75mlBtxTlQgNs8wXy6TDBrwkdhBAMA6TH4D
jSIDBtAJ1QWyDFJa4oh8qWaenlL9AIJJjSKhKr/6nAMJfyuUZTGIFFGRseNSISePAyhmKXW/1dQ4
Oks8fSddsldN2cWPBjpRjNqe6tcCBijnEcli8OYb30xlUM0UVMI+xLRgu4sP9ak/rMAUK2x1kHq/
rzo/bbIRuKdVMuOM12uVLssdYMYiPVYwDJFiXuf/4hiRHsQxHqDV7IDeD0D+ipyzypXzKwIk172L
T23KTfqxU5tg623LC/uXM3j3FAGWhiNA59QvxAPyAwb3CWc+zs1uQzfI8HsLosUEmi/W1RliSjsn
Jl80dpB3a26F8AI5AoffA2gu4V0NIVT4pbO58EOikKr45cFz9k5qEgEP2XrAkr18MSYtYA6geaFV
55biVVwIOnrerm0VBSGM7XRbotdXbFM3pfBcHpZI8JTd8e6n53fRv4nZpaa34MULEtksFICzz+It
age/PokCWRR/qzlxsw4vs+rOibzcSJ0E6l5ntGe8wxPEStG50wg693ue73qaJtedXZ2pVIe6znmj
RS5cz5jXYMWTzA0JOMaIKraI7gDTJxFRn7eTcZuU71OCaSZtzkoKccTtt8/TWQqfOc8sryIGDXPm
5OmyYNVnUwvus3U0HdP1ycwk8D+EB9ovwwp99BA2vbkBaD3HZw+Yi5ACaAo5oB6VhnMx7oNKDqSw
zX2PDiC8e+gxjB6d4a3WC2uSaSTbatmKcOyQa2mqC4FpDde9ae4/0iqqPTFFyh2vBZe3GZygqvL7
1goWER1Ep91iuzfBWL1rcDf1pKNdQZJ98U8u2vxBdL0k/Z7hFnphcv0Sj4IQSzliszonTW+8XjCy
ouX+iKEF3tlpOFJ9DoDzFyxS0/24azf6SYsiuSJuu2/R+sfpfYg/VDLxnpgefWHDPEQuKvyx5baU
UmNqw5r7tqhuHiELH3OZOHgjjjgm71fhLHaoYRswZCNIie4MfXB0I/S2gMAbMTnkmclGCJlpOjBq
9ULkHoa5G2U30oIWqsTV548xqVRpFDDHrIRVifgl9YYEGTgAWZH3MUop/FVmVd/Wz0SjWvVFSWx8
jmk6zxzweYQJIsPnEcRE9K0xSJd3oJwIlpMWJ48csDRYOi+J1UrFAIpNkDrahWgEc1GcSdRo4fzd
stcEHDeB3YgTHyhAYicz3xQSNGzrz2PhQNFHloCpS96T2yR6fhTf80nerfUX8zbvBhr8WkCT0Q72
Nq64qItkj/gixjWmpqhXMY80YxHjL43fO9E5L4y+EikiWexCKD+1qlv0gAH9l+kZ224j6xqUg/sI
9IxrrLKut91Nliwxn7IOHdnHiAPCaQ3BwGCqZ7z5tBXVRggtJVMhdydHTKbM2a9ywgD5ikgmWFWO
LeOxzR1rWUWo40cvORkfdqVFicPagfZyvdZ5UbOM5UfUpAyox8N5va2z1ZYQoF+zKb60I/sA0lIC
tMTVCS93imVNBuMp1FCiKumAcoBwtXt9217TQb5ZLB7eQPLjW+ICBoXLh5ewt/t2g7bUNRg5WNx1
VCOtMhgVYy0mUlszV2GhBFRduqM5hhPcCUDulwXIshW7XIYOPs0qokCIp1jP+isUigIb3sUED0nC
AnlGgb0Bxf1sIKkZ5A/BaWpr/QHXpc5M919LkeF+yw4CN6XrlVXZJeijnyphDZefuXVGQzCl5GhG
9Y/Nb0rMPVnDbwhhl8tZ5Cw2oNsn7lMTyigXmSxwSNSQpSZPrAWhPHDwx2cczCtfnNsXYaXGGzGV
dOEbJ0BtfuOjqiK65bTbYPGKjBnKQ2NxlnX/SuUqnGcs/hE4t4BprTR0aU815ys8GVks7t41krUK
U86040JZwbGNNaXuCPJJ+DdZju+3YWeT+VHP9RDwVSB4OjtmcjbIUKT1H1WF6fLp1i5SOSR4hKi6
XJR9ZJf+FTA0oZOvHWkB83ZXlb6E86Ti3jQ/H7NtylxgBGGtsXy8Vx6nnuPQ4odWyNfDkmc2NMl0
yBlzKxXlw6KnsQqh1wIXzjTvRWAdgPMCaiRUhhXXaZQZS4ESwcoT080n5eaMvr8K1SDFQbhTdYQ+
n5NLDlhMvAWsz0jEkMooTWFY+tEgXQMhJymfY4J4q8n+8ff8AKvs3zLppmWKNTxcqMtaWLGh6ZoR
xaoBIXSlXTEGoaNthiZBNJ32U8kHgGw77axIwga6yXTCoEORJ7KX9mP0F6Wz8uTHjKQxkuPwYFOM
9145FTDel7RZLKOM45sPS9+aHbgLTCWL65ncd/UC85hWydjWYyeJANTwN3KDJod5aVW2zC4/b3Mp
FYAGQMmPSaFVgUaTvylgVifXb7Z9TfhnbG6fPcD0eIGowlENtvz/Xnn/SN3+ONqz6bBzXtEyxe0/
JOZm68dNkPvAFlOmOCXQxog08FABcxKWjYpeoaGLK4ek/gSekDBiwRatKZa71vvQ3JmKMfEZhuCR
JejMZ0pDvLnpUf4yntgyg/5a7NHeUrHuRDdlJCGVDS5PDURIp6kaUtYjVoYxVnHcDphacUvqtzOA
Fkub7fK27jH4Tzcz4Bgcm3ueU+/DKbrtDCXw8wcbwCYpeSXKQRijFuQ4yluN5rhryZG72eXLaevW
LBXOAPFTx93+7MPYT4kgJZLS/tvMFK2yJDQKFsisrtDv8RphOMtKrHRJnj/xYk+DwGN60yESn1TI
CZhNfHrbgqSGQrMicDFTwKMOb4+Mew3othrr95Ebg/R9kM8Zfcg9aTQu/AMI08m3AE0X9MSMPdYA
HrfReb4xHMBsqEY6gn1x8HqjzJYuuM5qtrYEjD9re/mwezBiboPmVRdo7d7Rdj+KaTKGlu1xiVXB
KHm7y6sQftSIJyj98F2P6y+4arTDUm4qnXhfDgbhRHM7DoKrjSx1AoI/kx+xRiQOl3yquX1CwZx4
4FEAarumgkWWwdPkIb4O6N4J3Wyg4VnPvugzOoSx4awOMJnMuC+9q4u3Mun0SJeGLTShkJZHIaLR
FgouSdxOYVj6vluHNm++YbFU5G/6TXGnkkKSgkluVM812w5c++fZxzF0XZuywjksAjWhWxHn29EI
J4bYU/V8y+QpCpxTMPNYGkE+iTpbcQm/a1Q1sFxdAYL19mNA6qy+pAr2MXD991Y08lagI/D3vPb5
uyhFIyLm+xk+tzjD55UeZI/dRHNKbum/x5pozuWeCA9GVWW9r5dq1Ypzkuz21X2Do4OQSqR7PQhf
JKDE+K9ZdA0X5eilfMtlE04kh7NM7yCqNeuciIsEdGELIz/AFYoVmgbUcvrZeidgt938Irajwz2z
DmtFQwmsaCT0lg5QWw/V4P+V6upaJPlgAbZoFJnWPa7KsA0W1pxGbaIXtrSMvahBGrclQO6IwUgT
Jt4qTwiU60QUTZNcwS5nv6727XlSCO+XFEZHaYRaPOOihablLmr3CQfdllWClbIFppWqNSm2eZ/N
SqAelcNY2XTQrejON6bOl6AJgTQUCMG+0tEqsNIF+siYgfEY6W0oOGJPbdY4GOVCGTH+vtAmIGEb
P8TD91trUaLelFeihVxCwut3lC+J2svXc8Bge6/jyXYZMjenLDzUM60W7jQllvwgtcauSRa+fWO4
AZqw8DmyV19X5p1SgVoWXSluIMIzSzrCjHD0eUxMABg5qt/heTmJbWqZrkLniEJC39BhjlitWO6g
yE9TJReJJXLAeTQNtMRPsgYs1qm9tr4yO7LukrG2xCkiqD07uUtBlJ+RG8x42lNF46OhPX8mm8hP
sslnCzGvA1wbbfZw/UpsG08O5ktv7eCUeyFFclRjk8TdQANDPQKVX16Dk4I+FyxEtYZ3q+k9DkB3
2hG4LK2bKDsFyDujydK0dKw3cNAW/aBb12Q+bkF2BTYi3xEeku2IJa+UcZdY/CNvHHIJHMEjMlEn
PNRfxPM4Yzr/m8iQgm7s9KRTbCyB4lgQg5vUUFLMmWMguGdKwc0fw9FleeYWbFVjuAPptdkUGaDE
O/2IHgniNBKQvbLMwQFHbcMd29+coQogBMhtd3nL8l3CmAXmH1/hh2FXlnSWdQSoG1/Bk0VqWBHP
8Q7w4bZyVRaVTKmmc37tira7RGu+/jK2sK1F5UkyBOWjxuJCF2JLr6wZm4iAOk70ES0qE7mIxwoU
3bDSQ+I6LEqdi6Jc/TQ9Q/Z6uuM9rPQ7UhexEEDuZYChp2RMa13SFWE0N0KCBfoxZjm1LIrA6P78
eABspp9tIxdrOF3v3GYL8lw9cYil+8l2q3dwL7upWD10831SPfGIVRztELQuNXQEpDwDJIajF792
be9VrX7M1ensyW3mep2SSYLVzBodcizDLulBjtHMUYZs47WU3amFec9h5+F+F18UNn3xD97sx3ZO
MMQ3+zG3588zvVOjvcKuly5K/P7l76RL8mycH6S08efAeUePJlzP7oVEfCgS9LsWD4pAaPNEYRbs
LPVIKFGEmR1tDho7azX5Ax6NFQrsZbY8cwqpnXC3Ktzq2LWy2AEjzObme7dUvFudsK4bImjtwGNq
XMATZgc6Blqt5/04YZ3sZg4t+L+/FMI5FfIU8LOGrrEYDbGFcKOkx4a+T2P1pJgdnbuvDLed9q1T
CUVuz5CruWUu9hRf8NheydSCQ4b3z3iUJWz6/gzTw4zWjEuMytGCfgiV1/ypQHHjJC+dNZ8snyoA
oc+YoPcG0W3+m8zy/yB0lCkn5zFxUUY/qJs+zwriZPD+0HJGx5iAAXAjBY1K6MlJS/jqhj8eaVVd
lLoTHJjzgizIXVRaiykfm3E2NbmJsN+THoMIrtFTgIlSn5x+Nj+LnhJVnpPsUaSPeYycZ+jfS+vP
rYrvR7rcZG/NXNpt8tyRtkwu850N660fv5vXN9Ks++v4v8fYcLUVmN9YkF9qclYG9qmTNppycIwm
LUJZ4C5A+YQwoWduLA6KwMpUbmPZ8sxDlw6tCKuRhtY+JIdn+WgzaDEHKBxWCwQgDuy+BQG/UCV4
V1sgZ0AWZoAjjx3cfcDbdkULrv5OoHSQTIiQ44R2dZMNcazwzAH0lGJA2OiAP5D6i5u3EpzpSH/Q
9ynjkPkgIzm9DUFuQp92VQ27uUXZN8TfNVWZKKlumKUDgpDstfhuT8B9JqiTzrtenXSLzXECQqwE
OQPliJ3KVXOFEnhLj7G6BquY2pS5Iol6JEmeDr5EDROlon/hNOV2ARpXYdzveY62gUOoUx18FQLr
hELEQYCn5NbznNrpcxObYupFgISHQVAPy6tgB5vyPzCLVSxMbS1JIibz2GQMVn66XG1vsqTXr3nS
ypkPett8cEq0YQA3Q1+WyiMm0fWMbsJ+3BfCg4fwD4n8CgSlViGOxoAX5boJec+7FR5JsPTQE1Uk
qI+YHa48q08nfdVZOWmb///C1Bb+1un2DdOJP8qVFiHIPgOVuJnvJKNxRxBATSjVnITP+Qo7kOoR
8JXQtXoEfcpkEo3e7q5ar77X+q52HLcX948ydPROx5YOhTLx/wIv6yHNMK+tcpavixMsa/f6aAIc
nklSH4MdDLaB0liLVTKUEmzI3ftZ1JSQNmZWzgmpEO8PNWHVEKSJ8WG6rRb6Olfbnmw9a9kKigIP
p3NWcLYL6rP7EFiUqVTFrfxmWGFWOkvwbqC6mFG7BktKqX+6lPXvjbc5uHwNrPXp9HGcl1JZ5Ylz
ljbb33BIxGUz7KSdpEzfGWTOm/axeK5nUrrXxAzNHnTxaazgEQ2GuK0EbdDwvoVvTES191U+mMqi
dy02G8+XmCoqoDUj0LokM9JyiPzXm805DccDuy4qvVjIMN0TJrBWr4n5mg+P0qgemq0TJaAc6KR4
LhdlkzWsQi+frQdBKIsEWgg5LOJKpsCSTvdhEf8MWJtN3jXh6PERENnhPJy0hhWBLiyirYb+YUtv
mPu85ayubeYHQag+25sctVm1eRK2O5Ww0ONdjXKt0aapAsEMp/qaPQE4i4Yz6eiKcIch/fVIrTCV
pCyBstpPIQIjkNDxPKsrQCP+dA22O76ChmzcxJLyDQesN/2GSSgt85zAB/aYysL8Qo+AQTDLPahO
ojF2CD8OBTI8maBEkGzPSxTTEY3PO3W5ku+fbk6ELYCTsRfKXuepHpRZ7kQ5GHlg+X4jp8SlxP99
sVD3J+UocfmHApdqHOJOPc1VwugjaDE3AtdAGkHooSS1XViCQn6jNdpfEDUBVBQXs9TaOBkNUfm4
jDfhtIoZzJRiWD9vTfpFlXhaCJgg3TGwxJLXKK48CdlKNq4hsVUHJNjtFkNb/6G7vPTXTOLp/2zS
wy/jm9SKpRshjiizD4q8NdJ2yf6bLBlJKn38IZ2UWBZYkCTjdMc6TbiS4nht2er04ImqlrIMa6+I
RQ/HRlqWNHMHmMB/9Cuyc7yDVlLFcastK216ZtyrltB5bkmx21qoMqNgX4uB3SpwZOmH1Eo50q5O
9TPK2ZuxDIjRyr58kje1O+Uk5n6wq1BYfSbVY/2SZ2S7/9sXoOYu/v4Cy50/pxEYpGN/5N9TWa48
PIjUjyHQ/eZM/6J/ASTe47lT8Zq3WEsGLpBYK/oOjkkZ7kO/yDWcP3XxWueZAQPTucYqOQ/dZUD4
JOCOVYzr3dQXyPzy4aYTc7kQRagnFaO9AZIq+Za37/ahAB+dmvyMPM30qxfvYifUIPcyp3wyI4rX
Mmrx6xuSuL8nV8DXw/au5UY6/JpzhT8m853lSkpPY3ISzfLJQlxO82srqv2V1qfWg6nQX35L034K
1E16GI0uw4U4C/0mAEe1sA3RkwAReGSb0Xb+wXbWy7F3sfrDOmxeq3seyQTlMQPFxDgrRLCDdAKV
xxK9v4oPAaVVxwkkLLG1AEh7NmtVXbqOV6zbrTq1pRGpsvdc5rOCxcbppUwmmIG1pGaWcUPlvb8W
PVB0unspX9MZNk6lPKzFCFPvVREuFVnet9uUAFO/aSSdp2t5gIDpw3oc+lPWPJ2OtYiAWxP62YX7
qLEKHwjXHwHqOhSNtl89YmRk/hsJAoz3miFw0gcZcA1cWZvbZl3xIK1mLVuffwX/Y6ZJhnFk/x2v
1LHCimkyVYsDkIdfxEIzvvBWpiQVDKqB9usYlTh9s4OcRKIH7TyFgZ9CwfcI62j0oj5/Kemggn6z
0BDRHn0ePlSEJbyIIA+KOf9NF9kODw9mKWSg4vMNpUm+NCO/b1fdxsRvVqmzyZNWyQ1W/dnHtGR3
qZeKjjOa0PxmBW+rIB3bsJiYISn3zhjdpLGqDFzI2wqYuwtQl6I3RdSof+eJi9k1IkE1BhPNx9RW
blvNYTEJX8UBouapR5xcWGWr3PAOTRalhe5wzQwRXpbC2azwbQEGcGGahV7DpF4rW+392gtA3VnV
L39dDK+AqY/7puCDZ5h8s7gnp79RNcJLclg2Rg25Ap+hUggwUw4kV8Yt8AY4j4b8TE0V8CvvHGA9
udb3yqEy7x9qykabUOLZDC4HC8GM6ReMJodha/p2abl2QyTc4gWM3nGtSaYjZjn5K5twn2XZOZiq
zSQ3Ow6seO/UFqmLc+n+RvDnRb5aCeosgpyIZIMKLMW/UtY7KrlJxBivUAjnP36jjNNmf3eH7o/d
/UIaX3u2X8SH8cCSqUZswf4tW1QAOlVRlffuveDL/ZDtZwkYDBnfOe0hj01nHKHU9PZom2WIj3GL
jffLgLhlbl8x6HkHzyWZxnV7ao6QQLbcK/8brgD8rnuyRaEzTl7xLMj5Lokh2bUAX3qHv7tyHVO7
JsV+HX+bokttFASqjR8BP6JnGry1NhrmUc/nrzlfBIGh997Zkvk9R8RQEfSLYKu9tHEk3iciikIe
OLdcF/+0WAGyLM0feDI2SOKpoXvWJTaBE36ZxuctuxJaF6kPtkWRyGv5PxnHaTPqWvn+Xk8wuEsW
KJJXNBCKmiXzj55gWiutG7vx8FSuxMubI9cDe8W2dZe1k4fb8mfVlJuOT1+Lqc5eTerEzxiKD4h/
cO/MoyyEXso3tMi+S0FwFXMg+331MxfR5nOWO9/T+XjBzFRZ+C5o7DXtayvY9HpnbW0Zy05iszeP
/NGLnyBrauJOSBX1220wGdhhuczahzc48SZrgxojo0kxZKkNg99kac6Wf/UEp68pS54ln0xOuCWg
Yl2WsHiJkrc1S/vofR1wtJtwEVMabgoc6aUAQQh2sr8B81+Oc1T7D8Oox2sktyoKKlB5Jah+mG8l
BNwAcACtNzyGZO7JqfGebwlVbYPMfJ6TE0LNJsYYZhcP9nAMvlBJsb/tiJDMD6Db5zLBIj1qr6A5
VXUD1InvuLU+8WmWPmKHvSJ40RO5IEOqu1MO5LaBrqE68ykS7TdrrqBZgDTFoc5Sjvp63grrfkO1
hKSlQhKOk7gDOGd0DHfOHK0e7TpRiQNKjeWBeoEuVxOdi2+iYP+0zbfY88indylDC4mn8NVBNJ/c
cKNxDN+cpvi0LJKIM66cc6IuDjdMEA7WNbulAMyFXcEWesN9QaQ3Y6bjiiDliD6TZw9EOk9gRkpp
xyesnQVhL5H9jvWJ9bVVPw38mSjUVkG+chzqUwcHymirRaeRft78b1B+oZhqLAFOYUohHoFc7YHX
U6HCbIdv02xfifIWd96zDjKe67yyyg/hgmfuz0BLI11zW4FjiZ7UdsC4Zc6wMlIfN9EQap4kd9rQ
YR/LOXkOUnryomyuoYO+jzvuu+0rY1Qvfz6VqeA2Te3qYPBWw+CRZHwpnzL1LR8I+Dfy5PTse44J
Gn7EIMqZ8sl0KSzYjOzTw6go+0mIyub5Nk1rmHC0GaMX0MOT5vdUNiN9mylaNR0ygmDKk6czvtRL
NgrOd6V02MfQsry4FA6n7ENLlg6Dzl5Lo5KgOcyOoF9//6EY/vSqD5Ae9pT/faW0QKlvU8bisvk5
H+tDYKIaFcWg1fbtSpCx/Dj4mi2vEL21YMP9zxNi/5lDh+D9MmXsrwHxm/ZYzG7fzTMGolX9p4en
FgTvVQpmXD5ABDlmWKmQzW2Keg8nltfbu4M9YdWhEXku/jiZU8Mntva0xgeX7ia9BTUk711Qw+w2
4bXVcJqqgunJSiqZJEn3iF6imXuHW4dBsIrOoMk0htLA9Jih9dATSUtJZ5OR5NLljZ8iCgh+Vu1N
2lBjuyXvvSpkxIq42q304eEXgdqx6f31OK9bgJwr5kyIXKJBkMRYQOmXJC4hry56PZvqdl+ZmRFF
FNkytaP4wakWWRmTydI+A+JMbahbacIbQ2REufaQNQMHny79jbJyRr9aHImLP3Gl5r9x5urOeb5K
BGAQA4/A7J+SVSZu0aISF7RP/O+2X9Bd9vXJFg+qiMFy9vfM9LudLDR6Kqhls1iRhak7iZVPoSVR
AM9IPlMwkFRHLDwss9h9PYVxUdUPd572I0zKiUBb850PHL3d1VFip8jBcGxBW3AWvNbvdZqWCy2d
aTQCfTglRXbhHlQ0wD7IsM9uJETNEmo/bvv75ZmzLgX5ZOkqthAJNt+LbSIVnwJGfS9HdM0GU//s
5Sl6JRsQThV1CoPlAgdrlGOpKSIOY/AQXWV5TSy5/tWT+kg7iKd3P3l4g5xDx8yZXXjUuimJMLOm
573NdRsYQxck5bTFfghMBxE7rKAtzKVja/P4BOqhv1/tkHZaAZ3XGpW/a9KUlZQxC0Rbse+fGHQn
m4sSUauiqWqBigWTrm0nDIvqV+TELIHg7gTQgv3yxvHprLjbf4dhmROyrCDuW5H4UvrlrBG3h8Le
UrhowIJFpcGha4Ha1tm2Hjf7GBeKIE/lqSjPjAGraSlAfB99L7sCc+SjHmiclgfU4X8YWfKFpZjv
m2C6j7hUyCa0+Veqx0x5i93P2D2tE7IEWId1qWYV/SNYxBczNlMiVnkwRmUvQYk1B1W2P8kS2FXS
fDysWh6sujUzzXggNYwv6eKYYf/tppNUyRpOiKP/yTkNK4T8SYEgX3WkNUjwE6+Aa20g5jQnTe/k
y2HIftRks5Pa2YVWVoQ0K9qU2FX5qktr8NqPRr9lqQQtxFLi/qpCboEBBamfMhRA2SxGuYTfA1hP
K42IXLfWfWfluj6S1qvrdX7WBRHHkKxgQPpPb6407X0VdFDFCFjzjo27c9AJANNnslOaKEffHErI
fjDd1BdDWLdCokVFTLJ5iyWPASFZBbVEHbvQ5y2WI8ZLwaVOflb/fZNYqteLYhgBt/F13NbDCsFW
J69ED6GWU4zd7mHg7Dzs98SvpF9qxZejswfi0xl+60M5GVey27dMa5gequ//OvekP4h+rL8VA++s
graycHpA/KUbrFFHtGuHaRZXVDvdNw1lZLmp5aXRLAHVbdSWtYasOjlRNLsLx00WfpJSpOq6R9F9
G0qdUAiCipZtxUJVhpm76WYX5zJGAbM6dLtZj1StiaFScrT2yaA5a2a252x2Ev80gemIqQcfas9Z
1GGY/dxiAGMtKYmeIe9rSRWhQ9/lCleKC2syXRTUokzH79hSiakdEAaVys/EshQpHlElAHSeE2ar
1qh7DdC6M6ebPJM4h8IZBE1/l2IrSSEIEkeKpYB5bJwwDqOmgHDIgW3M7rNbpzrA0SpGqk8Z+kWA
KznDuf2Niut6/VMxF3pm1CShNaW1JDXiuga+S7QNMnxIAO08XmIhlquSgn/n+pPjZtm4QXLhr7XQ
Jsh5Eqj7WlfRhw+D0caDHbO5qQd/93SH13rcCXO5MY6FDELuJuQT8H0ScC0Ik5SBIvSdoN9oNcw3
4lkaY9oRoYvv53wd4WKgWlZ2dIq9ZIPUQbZbZOx5dCqh5lJHeQMC3cnPT2TFdgdO3/ZeSfBc8vNT
46FuJrtDQREQQFF9XJWNRXP4AMrDZ2JLo3oameIQEdi+nA+sGFXDLkV4zCXbMH8vJ+nPQDt/nfiO
CXry/BF7PKlveb6m4QST5yFnaaENvdlxYojd1TKAfNGezarHFyORWP2OHwCSbZcLxAvVUAGwUK//
dvWfkbBMjE6agRspaa9Tzo6pGwTMlU9tJM5jjF1ExhqEu5VtAtSIrY6/+NugD5BSpQ+sDAhDzbbD
FpPJ5aTdTI8jn+gMFKYoYXWsG0BanzjvYp5CLiJa7xzdTkBhhDwtmrm025BkODvZ1kdl9T/GucLO
IvATA9RJNXnnPhr5et1wku4pjTpLggof81VO2Je8gibL67nfnZtmPVn/7TiQJcLd1JlhEQUiQKuY
1Zk+Vjb5Ix6ItTUZxXlknKS9o/r85b60FKko7qb2ATehzEGFM7yB5FgjE3yk4T7ZTq8EKSAAgJoV
VJTMNI3dnqVckxP+c5Ibxeir2nGGx/ytkMw6q0h7B8PPtC6clIrBVABvy8VMcZZZ8Sn3ijR9e3yi
UQuZTaHNyRIIvGkv34Kb0FTeQH8kFEQRnDHs6VBA6Q5MByRr5d7cry3o/hASPhQt3BQbhaAjkPzZ
aaySL04pdgB/9HUwdAsBGk48T3A79RHQxSNsg50XgWH9HEflknrbsti6XXvqRVHTv4q3/BjIhvPl
sEe8mQIwz8niV/ZKQ/5UHjmNWhmAPFU7FCMyn856vgj4/CWmNDoBixzY4Lp7trNXCuTuMcr/2Vfi
Ct5Ew7UTF6bR7K/Dw5PuPspNO2GY5EYJ6QGdyTCLbwfEwFliwc92j8x1zN8YDPklWqqP0I9cyibj
1JzjWAvATvow0OvpHc1TorjLKIlDLkyDYQo2SYeGIopbgbnOoo9Srn9wH871KvMddY3xGJ9bLuuj
RfP2D/9BdL5UVJlP5YA2awlkcbV+DBcZWxujR48PttJPyjl/miXwDalfLPkH0MQ1ZS7PxSQy9v5Z
yhXDxL7RtDpwRG/ymf2VWB2xqTZlQz+nBMGMuJVbrdc1oNTYk8fJ/Yoh4VTKksN3kgFqi2MbDywj
RVZRWuEwG3urSz/XtmjX4czxKAOAYlT41SRSRL7Fi37ZQjVIsCB8j0Gi6PtMVyH67Vy0tbmr+T+1
u9IqQYhyiejT8UavGJzTJKsHPOKG6JUXEx2NoOmQ5/AyCBFjmxVIqXn4KK7mclzQJbFvJo4gKrCk
jUmPObQOBOf1Z3DO/gyYYs+kIfvWfQmUAwSmaSf6V6EYNZgGPJjvZ3adymWhlYt573V89+VvYNxd
dJFItj/Mzgtyktcb0xlzv8SBsVWBbimpAB22mbR1WsvZIVa7W7GktoYpSxoPxhiOqn7m66rwFqdq
oPuYDlihoWZ6KI9ZPUqjsPWkOETATC+xESuLr+oemKMZl7ovG5fL7ApWhumwL4NNU/DtQzlx2fUO
e0s8sEPRvsiDauDj3AfcqZmRQgy2uM3ujj4yzXmJCtz9RkwBdYMIM2I3RThkc5Syed4sZJLYEgxx
3eKVrmTNyGTQJCS5dN0qBwf5LCdFPzQqt0z8zu/j5SYnROWxTOmScvmrIO56jQPE/E0SQAzVHq6Q
gKF38kUWChaGFAfwfj/VWamOVQ92nbHzIAjvQRHAK+2usy9uc61l6BnmCooozVuRFBiMhyZEAiPF
qg3TUpVU5Vl+x+CUczPcsSCOO4QUziH9c6Dsad+X7iXePG/ZgGfN+UwDjvOmbRQHK0kz8ytawl4Y
EbMZoEzPJtvYiLsU8mnPQJ45zyVpJqQeFAAXejBZRQu/4dFuUSNjr93/5xbdbC9DTi5ke6sMUjxF
+ix7lo/RBFVZx1FJvQSGbgazXcProVC5BN7GzqWHPUcAocILyFVl1JQzt+SQcBxHUxvFacc64lHT
ewlbKtwhD1n1zeGaZflpcHV8DNU954aTS++vEaAccrPjVcYnBarOGOcV94YOeighJgRk1mFIW1PX
8KC26N3pIWEJUbngEuTZRyROsRE9FcDJ0FkNvrhhmYqLXF4nPaEOThlywe8ljv0/bA1oH79EWaMe
/u6Od2W36NBvkmCM4fiE/SYD1DM8jCKPkql8y89ajTZrYX3RtgW1iSAoMKBDcIlD8nVEl1aDyFhO
WhFL2N045d836idy61hrs4uzQjN8Y6flhGofaFyM+vYfqesrdJooavOV/1qewFZRI12WbFaS184s
LGRFyQ0HlK5Y2N+i7jbZpfeqYJJJ3e1vvx4XsYd+BYeg5k9TXrH7I+QiSpenAtPBmMcvrBULJond
JtCokByORzKCF4yUQxX2p1GZaFGx/+UkedpG4ea2fHOKQNPB2xWYjyMyJGJO+QWOW8fyD9vif6HV
IeDJY9CpHZbsU5AKu3INbuAkcSpz5XJTqS0Eyv5cMwFcXMVR2mqsHPPZ3OZcdD1nRD7KWu7OaKUI
xFZtwtw7hnHLkYtG6enT0FP4SR7oWBbzVuTOKiq53DeRqOjyX3OQqi/c7FdrG9yY3M/XC1jpixLt
EsLvJORneDe5JkxinF0K0wRodK3MGDH07+ksjvUoY+oqyS73vxkPfwHzhxQTLU+lsgGwIulXLuZd
ZSRu3rT88u6+wdg75ZFS0EdMHN/8575M1Sb7X9QURG/66ihbZMJiiSxsVFjzaFcHgYU4VdZwn6Hi
2fAze7398xOYMhFMmHGKc+4T7WQ1OE3brUTTYjW6n5wrzIdj3G4u2FQkN+tcbPk5JyoaSyhj/m9X
O98uPZjKj2L7TBD4lWXs6gfSxfLgBfw4D5BWfbLc2Xx5GDwNAiMogu6BQVqvoO/8AKNF9JTG7sYy
QVkmqsQyq8UbuemX5fMIugiDQa8BsGWMW2IfywC75PtpSjFbCZEwU6ud/SrNypaxClJzD+ezQcQ6
1jynAItAUnGPjWWRn/wemj0/buFDa507TMRhmTU2PQZz+6e9lnFJRX0UNtSoRa/W7eqtfQuclg+T
jVkX3i+b/ddVNOuc26SWQBJpVVglK544BqaE53FUZRDGwGzp4F7fvjGAHJaBnTFgx29MAPQs61oS
IUUtDTfeRvPXY2uItjLA751B1j4qrTExhp9b5VLZ1C3S2clmlb9OJMQFCu/gse9/ttea+Y7a9YWP
Zu5ZyaO57uUvTJrol3ZzgLfjdqMrLRLmV5HemuVv1Xj3lSU1ZMUkhIcmvG9CDnI1Y7A8/EE3CDk+
V74JSupO8ATo/7vLSeVg2PTxls4y50zkqDwjtqwESeVprvJZGtzZVBwuv1cqUfgteaEQNxBba3kn
JwKznKALRzCCfcBEk5hhG68SpBSif7v2oRM/yJVGZntD0sQPMxVE/j5WMgMMkS/duj1MF1SA+2Vm
/4HPlmGy8rTM/KnqPNKJ5RO0faP4XY6/fZ2JGe1vILOQWC2tiUlMq9QvJF9j+b81HwWXggqUi/bR
J2YuXTn8hwdE5MDAJ6BG/bSrkIn60mlC9rhXQhpKpGz1P22YSn61l1RVNtTqfQXcvzDMlMHIyoMH
H5iel4LvLFCPGbYCbbiuAYPSvdaGqz/hcSv8gr0WmzM7DghWPC1JOva3FV/m4ua+dc6V9KW4WKw6
EF4qrKIyiMNG6x9AmdltJ2qVB1938xt2fXtYsoblgB+CaLivM2fYKORbq0D/VhkPdeI/3f6L3iDS
WinNt1/1xHPhQhQCrjbRwtg7hz6zIbxw94kB+8ekQZfTt65QkCVmzCAawVpI8JkCS1FYd6tQhCWm
Dp/11UFM4TOxXP9XzcHJTI/hxCQ7kakTcPg3RXjTDEHHFmsFEuMcpJrh5habcmmei6ymIHqhiX4X
BbdtOer/bLaIkkJk1EJmSK8Tlq6Qs0RdEh6rA7GIM9kZKEgs6HjiVTst7+WM+QY6llFaLg5BJQnf
NX4fv+hmx0BTfZLGmAzm3rFesFgehf0M5ozDg05w2bxeLnY1NCBOQv7w48VJ+/Peuj7l1he3tdWE
iMhDSZtXNTe54OuM5tQRCancRvpifjNxSPbsEbnk9JLfdWYbSMyKy1cnXRBcQa9mNrHwDJ6JazGg
fwC6KYsH88WyuD90EIHSUoCD6clD0CbzaGV0vVPuPf+Q0JDcSHVHl1FLu08A6cDNQuBiFcU+IHAD
bb8o6kn0nJ3QMeEHY+4hxplzzncbdqopdC82cymdCE7UQfdjLC8CAbtOJ8e8jr0WN50nARo+eDbt
s6WOa0SYfBu9XQo32lTPBqJGWf1ylkP336l+VJ04nj1HxGB0Cvf20HpT6OwHK3JvdyUTaYh9Vc14
kDy7Jg8Zz8a6+pye7RAycuvxsyVy6VyCJeN4Mv4NgWyUCjf3X3BeM+2YzM7yD/0X2aD85u9R7Mvm
jHJoXR38gyCJnFDJnhHZAFq+vEcbQVb6i9LzOyXDcPJeApY7foIhjWqIQ+ZtbQPkBGPBz1VhQf9Z
GiUPYvl0NVMs+kPOL5uUNAjNYXawYdcYJroqIc2kBgXPaYJ/B4lUx4S9wtkiAvjVzSMd9wRPYgeY
DBR6a6RPJ6rbRcFx+jZBnk3V437SI0PSV89cncqhJrTff81VCLGAKXFfWMPfj9BKNMpXYZ2XPOy/
l+nAck9npgL5PWHf6qOExns3iuuQ2cNlRBJRbGR6htaaFjwyKRfNj+TrUjDbjj/SPY6QKCyfOVhe
UVAduhJEwNu1UnacBwUgtgTDzpO70LU6kFjE545RMjDZ+9GMxBHvdKjEbSSMCbmj4CFuRCnMyrri
LyiQDoFpGOc+V/uFr+5Z52Z3aGAr4pAcG164QLR25hjAVS2+DIGobbNJ2g5mcrQbxKbRHllLovsG
FhQNzitaOeox1vC6wdn2xdU2JAl0D3HovKLbgZsRXdscAlWeydowqKeYYTVwvOybdh+8V1Jt1yf+
QtWrFNQMtoBzbn9AsoBhXPzVtAZKJPeO98PphJetbW5sBhMs2YXj6XYcEhxRYBFYnusZukhoCNPD
lKZShOZfucPG3/TvC2IbDyJ9zRDHm3/B0o4mQMJGyN8qd6QrFKSTGDmFs4vHZVjfu5s6QsxCQEth
WK0QvKOSCJs2KGewVh3CAhdnznn+YSfvoaNwQniiGRG/wQyqGpEwmDKmSJhUqY3DAYzFFM9O3GIe
j6PUAV5jBesB3oBHgu19/Hy2Yj4DZcgEgHloqOIwJAr4n/ZOWAG0MQkTA3rMJetqO2P7SaC7n0tb
CAvHglYL77c84rX7Q20yzUQPuM8KXEOe3z1YpeKmrzkKFoRYqnZYIvQpVJy3/ZMR3C24X2Qu+UxT
t7PZJTtpilccB3LJVF4ULdv77wWjSTCmnhKlib+ojF7iglC+z+4/WP6Dp1n5E818KhB9kaQBDsg1
+PMP/NMa0aC/30g03/GZXBv55bFaEccMbsyOlMcqap0W9l/JNWOwBel0KJKZXrTAvcRZQnshzCLZ
RliHXEnabOq7M4Eh8SAUiRL0QvUWGLDtaTiLHoCYv+eGpkxhVyVxzSn1SLDVT3Z+dyZcU7Ta9TnG
MSvKO0TSrDxGQOmmlZlZ6P0W3fPp9EV82z76Q8psvD5uiz9zf7rYBOIRAMzC0K3LRCzBLIWk9p+G
R0ZI0Xw4vICf6mmZS0ULonwMdNjPf0nCfIL7HKlaIXNMopaG2Nb8ukoDthr5nxiV2j0M2Evjz4xq
MZgBliIt88O0Q5q1N9vsqwOfU6CwJkQw0irXzDOnf4/YwchYW+3HmF/DatBh96nElqWVsCfIslvq
Ao5NzYrlOHDb9Q6OQ8i0rO6egpngjGJmVruSndmg7TKRJemzq8pJFEkS1B3QNU7yQUJFFU/D7OcE
xvCK2jiYxFEMBAeO72hy6AbwJ0KgcRpA5vjjn/gAOLzzIbyONfGnQ5KP0iXDPR27s2y0US6GSh9e
Q6fWh+c86Xv/zrhvKd+C0SXBD6XlUxUVHNuArLT0zg4B1jaVrdfCxp2mqspUrV2tN5ERwQITZDfb
8hAShv1AwswgDn8ly2Xyk6bbSYYFaSUKxRQiX7LVzHJYIuqzpNAVe5Pw+kjEznRMA6fOiDUlfg56
R1EPbeyOGHCh71p+xJ0hkQoWLJdSWwEbUjUjCZYdlTaNpezs9Ip8FLQxTg2AnzeXwPM79bS4BHKa
rgBEcqD7H/XCavVwOx5m2vmFxfyTXmg2VVwE5Y02yPfF7yL9fws4QIpccChBX2j5c04Ct7X7C65A
hHAszmpIA26Trvg5IBbPbtV0sdOIdFs0G+4mXnF4ckpFYOYut6lHys1lufkCeYFFA0FrkaghR3mh
JX1JttBsWG4R1/6iea7nXZpxFViRdPB9yEt0FW0rPSAqe3exMWk5Vh5XoXK4phC1R1rwcEiZJUzn
xstgzmQ+c7Ktlk2ozGaSgx30qyDnh4TlckzNecseyV8DaeAfoD+OPOKZMaofzEWapukRPb8T1oso
QOkp7yzEiQIK7ZT8ZFZlq7PQsze/AZ5ovQ3A9I7OUIsiS02vC9ELKy5GDa19vvGQSoZciz5GdIMx
ryCLy5fjt98h7lY3I1+CiLH+CxAdIML+etY3M7grX58dWWdM+MJ3gYqBPvYKjvB7Kh+nHaW8aaeh
jn8H9TKRxPyBAAcCUZbIJjDm73/wSDIBMafCIaU5HTrGZM38SwWV0A0K4fp5KFHnhVqSdomenoe9
HuoMoiTHKM1WAzECrAA8NpeV+h5ddnSIANSgANpDermuCyGDeA0QHyR+Sxt07MQvrXSj7g9VxaKf
fP6IN3eUg5AjQ2hCyQT76kxl1rYHAl92ssONSo5QZ2iHJ1cBOWqlOo77pmYSGFTOpyNunbpeJAU5
zl364AfxRFDlAzNIpSZx6HzbZ+ekUyLouujUWtHMxEQs/e5gRYDGJLn4L73wNNWzX4UQ4xSTtVD6
lfFrwpv9sTmZ0ZoS+ePb4nnsxqSZ67RGRSRjvsSV7cqcTfD3U38dKZ0Uf9aHVPPyoAJhhaRo8FYx
MRC3PIvIFk304OgqgVEV4JgsvF1PC+4DbzkqCTiT0+Qvsi+EuwjJu6vDlYB5bWPVRWQzEv9ieymA
0BlDig0N6T311mJEeTkgwN2UOwphVi+DQgHvnm5vsD1THD98jOyxapZ11sgqR/UQY+xnFUgRPdzd
CMaxJV7gABVZ/XoV9frOS6kd47HsSImNn9LF9cl+kWyGATmqgOWsZ7XswL0m/xH9JV+zZIBnP6Oy
UeBKdg0pGQylmZTTREoczrh6DPdg9yqyUuf/zIiru4KTPg3rsvMrrooEf0Lm99MQwlCp2PmUnNTB
0mKjlkmVU0QA6nL1Nr26MsZd8UNVffaJ7my6nxm/yJsfX2iCTilZOU77OkOZZzq2OErEJtUJ+2Tu
+D57W348bUCqs+vyqgmlNkXJ5YHLdTb5wvpG6w43fT7Uofpy/aTOt9xITJLg6awFdwtQ7zA93aeH
wd3wN+eJvQNhuXC0nBeddX4p3nVFM6696uKcSFNb7Pv3VpMLgG2JSwqoVyr5deXAz/66KiuYaSZC
87SZ6LxD0ifwiGoDUp8Afat2kk0zOUoQVWSrw93ZJvaUeJ6CeveuHMyHg5RpF06kqZfZyj8O4P1B
qduYF4vNJEDd3rkLjZE1JAwgRTBD2ea9AuxyLAK53Un03z3RyItjbTH5TXamB9qYWxcQdBxUYXks
yIVYNKut0+BrvSEGOYIJLXzC6GPLE5HBrMhAx7gO9Lcrm1tLQamdZin17Sl672JEK9oOTjF2fFtI
VB6VruvF6RxwRlFahAMNbD3RTCFlIdR4swbha14hkhF669nDQb7XfEQ6MLRz1JVLxRNgwN3hlHb8
BX6Lsvl4kRJcmTXUZeSX0cK4rg9V+xIj5I+Lxu9a9Tc7Smr8Cwgfx7EC2ZEpnxlGfWlO21WavdA2
dRskdchyGZbJv7e/AqQmTvDWKnH2hDjUsqQOA2AWZqLq59chFtOwl2O83BWGoN5hwmboc1FpnS8g
XbevhhKYNEuHTVaoXw3tlFtDBnkfD2oa6FF8Anf6hDck8IjATF6H8UGA8CFfWPfF5OZuGNNxLwQs
Q7P+R8VG8XomY+bk13jR3k2IKN0JcQpcto148JPxf0Hake7kqw5Y2ut00Raxh1R9hhmWkjkCmm1S
Cb0YNRUkmCUWGU7toOJEUmNjGIfHe7DgwEMSkk1+kcZphF4hrIeYMrnEYpdhC7qQkBfDuXdF4UhU
lNGy+7OyzEM9mznNX3qopqarTkyKdXDtwtF1wFyalEjWfHQwARrGlogVBR3lMrnaKa+Az+uFdTKq
ynN+K4SCwm7RJRymPMehlE40KneVQpn9oOaLRTDP1ZG2A8R1frSjelhjWcPzhYHIwtPlVLuOGp4c
tjsZlrYSBatgElOJ4BbyRbjmiY3tSqHIpZ+R9lq8M9OkhrIiE5Zt8HxbQsJx64rRHDA4nMP6pA2S
Bhm43gzhbRNauKZJZboe0NnNSL1VFHDf/mLxfpERwsVU15mnl38IuKrPqUG6sQOkeRIzEGg1WMQk
QtJoub3lQzF4QlIPXK+mIXTQxrrJIRxNi7rBAC1me49zmwCJRN+u49RmXMs5nyS1g+nnN/k6B8U5
LAzf0p0sraH/ONlWgSP9QWCuhOqXGVb8QPt/n7BPotsf9CjA46KE8499RhBiy+1SPnmZw8d70wgv
sy1VjIeWixfsj3MwJoM+skSOSHbdFdKzxsCWUjMTV6RLR3slcBVFtOCaYEKbzOHnWF6BteMogk3e
azd0U/aCKq/pd+kNSV1wvcmYYJwlYfyE/LwGuiqllA+k4ddIyZ6gaqjsXYsCCc6bnD5e0aB+tknu
vfx8iGMkcT/hFlBxfoKQ8ivOMLRDWaF5/RkYwvHsdHA8Ti+99P1M7VJIphJQk9QuYuF3a7MvidNA
xJVW5cYz5CLatOlauLn2qAZWr+R5LNFcv6EWzuh4hxPlWLM+6Vzg71rKxGn8y0/DClOnAJsc7xQM
hYcKmvsLW2ZNGotw2mpXWUvApVVFivSEWVkXnPvEqHgUT+tCStiO07PenwDmz2B5zRD9NIeU4phh
5SbuDzSEiL6utMHSiF/uLXRhy0ZmTx5N0rWMiFwVeMfcR5Ud25i+pyf3ygGmtmmYkAVe5PbfbUVF
w22Xh9JmUkR4d0w6XfYzlEic79640rtviyqlujQmpGsfqDehK921lRKWCK+nb8v/fNl6hJrUgv1l
bb/7dJJIJiYODAi9CrDv61vts1yWDyDznlQ+k2og+GnQpslRcRJDSYYrKIdKCSDCDCmNZJLFomAK
EmyNtHwqjitHApFD7U7xp+fqye5xobca0QWjaUI/pv1W5YBkVHRrgpLATD+rUaC7v4bVZeQW9OJG
zenxtFG6l+6l+GDIuQelnoKgxI7dJ8RUp8hnINIqsww4Ho7BUEl+xW+EBcMRxf/GARv6/M12y3+s
/WJGGwZws85Cm1xDhrscyQNzA+t9TDDxRUnnMOfpxF/OSTIP4EjRKAyozjWERBk027PCsSUbbCiE
AAMi6Qxz0z6Gd9i/eBOzVBuSmN0xUwHRX3NpBkaaNEtbSgXWeBPP1HS0hA9MZ7j1RASpCu6oWWcE
sHgMlFj1b5Giu12in3cpSIn10rHoaQFxAgj/2L+sLY7rhmxzV8I4j9mQfZypiHk2vrVjpoHucWqW
dmpr+l5gtCW8SR2nRraQzY8aGYyiTk19MknnBQ/1gSg6WRRuJmt6LtoD2LJIRnx+2JX2jeAggBIw
ypFdk7cdPGYwjxB5DE/73C+pWTFhnejHII+ftCHLYbxwZ10h+pNRssykADG4yVLqLKQ90+SxlOE/
ifFoPLZ2SylcQMKi2mM0JREgA0Q9gKWBeYjOLXe3QizpAKMS4v8K/12AhiQ7rQwT73CBiQvMFHsD
EIPtuE7311jPZ311BXCjUJlUA4r863XymFjqhD6/dVDo528nFWneEub0jnVLy7t5l8Ag0fSoKGmY
0oXiGCKettMwAuLgu7VZ/l4YisP9j7GvDJKn6Vyg7Ua/P5OVxY1gchGkWHtLRAJXrcMEepF0u4db
kXiXZMj+QWukLw2b05YrLCh31IugwSGPKQkeUnmMtn9mKiJ/GvBuPyBeoDK7rSEXcLWq5DRkH7Gt
JQiEwn1Ph/IauH7oCt5bUQtG7vYmBmLrJlwmJk6KX1upbAWP4nncN0O7rFANvDe4TZ22vCdh0DKE
I0CqaVbvUjU+fueATbMNeDfhZebXsORgbXHdDnOKlFJZhQnD24TE4XftgOup9ZegUn0q19Z20LBz
XKoMaPyGP05v5l6rMIHP+aPYKOn9wsniL5CM6J6AD0vABFoJUZOlkfy0gluVosqRJ6e7Q2GcHAzh
GmVCtI1Z33SoNUZ5MyCrYspNfjhbtQqYHBc22516rpkbThjPj4Q44yYY2Ut5oH4NhzYU1I+xQQtJ
3A/+TwWHBc1198nH8prB9/FyJi4GnP7c1Es2PhEE3hSHf7KLbGanKbL/JxRg/xBvA4d+VSjcIpvH
FdT75FWenkc/7CINJjkeW+YNrcZIQIieCM42MTS1TNTh4R1JQURManNH/YsLrNk1UqkblvPamwBE
gxoZ6Oc/dQFHS9V3x8ZsKb4zhnCB19JT8hD1/LABIybwctwSCp6rUcYCsyfpeIPvMCftIYHKMr1c
06/SqoUrlOOKVNEhn8JuhDleUgBMwQSZOAXzc2QDUHzmFMJ2jd8GF10dEvMzpGIz+DbdPFQ4r9vy
G2FY7GLDEAzAZSIHFAR8Qqzng2jbyPthvpUpUyMTzYrIY7YC5IK7Dn4bHb/UIP4zDLM1hxXCelZM
vkGL6yu0X5IHwrTef4MXkFiIZcV6kjMNZz53mAbgl+0Xc88R2pzXtZ2Mz5rCg26id4XRZSKmdmir
bzXUjq1Re/3FMmY8rFoDC752yLZYE7NwED6s1GC5KLj5nrOJSR4Fvhdy4zWj3LQcaDPgB2A+bH8G
nwDbb5/5IDk6L/RJPKu/GF9b155hcmjg0oq889xACtqvwcT+4mu1fjV4lonmliJQomObCL8BXSuv
l08cnQEBpH+UXLwHDum1Q+oQO79taZ7nhNmL1IspfMZrWHzIQAkOKl3r2dkYsx7GJwJ+QMiwn4th
p5YnZdK/j69EbBo0amuTWub5Pu3hTX5E/qpPdE+JTjK/tkCnyE8JwNYL1eu1OPWnkJnsZ8ivCmQY
yujtwWRZUOIxLKEOjvrnuR/X6Uw6TN0ebWPR++0hs0ypB6tDfFIka302rOeMNu7wqP4Kq2ICpWPq
R1kEIXNBd49C0jNXHf2k6aj2YuC4guW3Z7tiezDgVnQtwIc2CLIzipOehbLDSE8HNfoB2d1mKvun
9+AaSlM7E2i3l+ltdtc5hsEvSweVcpoUb4/jLQwH4LtzvdfyDGhoN5IMVTffPoR1wrp9cCkZ5VAu
9O6oVPMemgwSgnyKxURjnTVBjjZSjzvx+BQMPL1IpCS2BXlqo6ySVfGL4pOaeGXe+xoCt27ECMvW
6lJ4b+nS1sa720tAYYz229CpR//rlP60qdRibMVN87hp3JZBhJekt85U/7HLre7EeaLW3iogGVfW
yJ95q/rrTfJMYlOt6nSScAMekqYMnAgPm8zK2452afdAz6wglmmcEEOLx9iKiR1njaHnroZ95/Co
d5OA0416G9jPMW7fHNtxjxRUdyqVRvqaFhGGXTOfTYVAs7OWE5QeIOCAIdNMK6p1vgbqcQEtSjNd
jnzuokXKjYrEORZCsaAmJblQ8PNRamW1SmmNCPqPMXtUjJqBEZKpvZZIXJhCx/lJdLabjOVo2FL/
BffzNnfFqtZ7HzE60cgshoAe11FPPiaMohIG4FJ7kujbOxsvYeWqzXXelgMVJxYHuDqbbdh5WE7R
ntnMaQec3Ne48UHyLtUl+henjvfg4rUpQ4fmEYryq95C85Z5fw2ZrcrsEJWwqKN3xfYOuoS8kDLg
8Qm5PUKuX8yEtUtVkyk8jTGIQ3Cn1T/m46+uFY0/yLTXQEjGNf9SsJ1Joyez9+RB7NyBYIgyihcl
qcQIJNNLa1HbNj0z0YJlEZa9hnIVbq3o8NJHnF+Zc5SVDZWGiw8cGSfW/DA3HLzgNi+JSyu2p8OJ
yMgYK57AbJUrDScJ3zUb6MDnX9CaoW8Im1Y+Rjk/khQqtSODUhbx9ORNVuo0YHVoZAAvb59JSPYD
b1wF72AIYUQMQzRRvIU4g7B14/4ddmNeTdjFInEVyJXh+5q102V8EOqP2ZlB814/JVrTVIdPO4SV
wBbTfcCbOnJtpz4GJbwk1ArOHI4ooxlVIOEerxr1ENTx+PIv4MruDKKAJIAXwDNaqLSCFMocMGq+
yrk8SHkFnoJ9DDZ2KV8340c+yeBo7fX9l3j5pC0eTIHJ1dtrvUqMC+dDTeNaRSdjdSe4uh/qFDFm
/R98PqqYf1JkouYPcM3kkDnM5QBO+p47w4AaBo1XxC83TOP6Y2iS0PkifcJEXqCvoOuDuoI/+iex
swDaVcNJYHocyPpnxJFFuGR6L/rO/cvfOj1RlFOCM+g6Q3ZSps0C1gGJ+3vUO9KW1wQ+7tZD2NMF
aHWgkNO2G6jhYwoAtXputs5QGbd7IKCHqkpOzmJuFrbQpjpxvvBXCxUDxa7veb482UAjwD/kXmw+
w+B2JEhw3k4c0Xry0WQGd1olg4v1ZYRUtH2+JnKqTOZkPPtrwjGAWw21kuc0+r9igJbTaEkpOqut
Gegi1/PS+yzEo1iKjBnfoJYubYdIcLfuObYcq45zJTSWVyxttnK5HQpb4iHhfPvXjexiuGDfcB94
JO6jgb62ZL+slezvrUJqjwyxW1ZwwT7tJzFElT9OhC6pOYEFfi1QFSko/c8kpAi4siTd04GZDZ/f
LhSx/b9ulUnCRl0NsVt8eL0xlIcb/ndryYKk8hLj3iColG9Tg4tqAFBeCG2ckdSF72V8vRo3z6vh
MCaTUOsGnHoYhvyvnfypZnP3AKKl62qdjpfumYQVKghw+kUObz5TqAQ5CJ1/zWibqI5uGA7wNaqE
SbNCYlObZ6R9I19gNDDvFRE6L1Wwnb1Uk3u9XWGis38Rb8EMGeCbPmsMb8UbyJBzgsW67Pw84A00
8aXArqFxvUrOHt41RBvHP+kabYUaYIWsFNMMhkLwLrgZBMoPkboa2nZFPbH2OTAHO2q1AyW7y1pO
o7Ob9WPIyY7zTI5WGsLAtZPK+N/5KOfzBULwhywWHWqyPGhus5TIWYMwNbOsHKxFSiJFxBxmp8Dy
/pEv5L3/hbhpnnZxEN2Mrv4NwnzO3/UU8Qinoyl9jH5+WSOufvXVV3zd73rdZOWR0pIFNQeb2XVA
TpC0MaTBoRf+Gf11E6ukfdY90Qz/mupC4Fne0gKeRIpbaADnuCsK7A/zjONZ2B/UTLY+6gTcXleo
GfdO9Zzbumzb+xAMHJLxdUGkePCTS6gz0ojnl9gkl26vEeRZpfVdAcbe1hnrHCQzM+ucQd/FCEeZ
40XtAGKix/nccMf7BfS5H46POIy2cfhkZ0UTKdlxOiWSJFGtjdwGTaEPeIHKSGUNAENo+kj9OZEn
zoCjC8tQHPLMhXiZPLqy0ho/GPNxcLgztoNQQQJ2wr2kVoU33tyHo1eoZm/F11+kCnzu6fwM5hfk
4IazLuTiXUXYMSTPMe/Xnm67+lKcoF7eyoLElO55POlBRqyv/Sbx83LF5yAStomVPiAoO5vqzoHJ
/Uu/JQHJ9zrM0RLrRM5bEUqVR4Hq4/K2SVDPVgtwGilq29RnUIhJ37y1XVcHvlmY5PY2tGRO7dmC
0IU8V56MtkCcyFTATfJM69UD0uYgdhfqVHhIdaPC+x04XMbfP4cLITKkcYirfjyif3iHFH5vxv0n
1OKUnd2GjGZPxJfH4viFXO18nq84He0KEosLV2wzSIiXGKlG8FLrv3aZO/H3v0o/8WCcmIM2vmwC
QGP15S54dI86Mz85YX18aKbCLBHqATZL0ikfaPzJSGRF6iMNxN5hQb3TY+arvl2bbIWKrbfeXCEo
2Qm7Ite3L1xNdff4Az/oheX63vtBXJ0CL+TX0n4Yt/BHWWRzRB3WliZeORCZUI81WBveqQV72M6k
/PGC19BElK9fUsAd02yMXPh2H6T3fDLpJXsM0AZUkaW43XTRhz4kVvWipc8l6JiR+IeWyhrkgGFh
QPK2zbd0OtBOT7CKnCHhcIOBoP0WDekM21gBMh3WwshObvyRb/0V2gDPrGhLBubE5M4qL/ct0oDA
bRZ2DJB2sdvHFO8n/hzGYE+tu4n48TT1z8G8mSLBq1fO0Y76iRxowJ6hIMakH6fnGtZjJm9hgiBZ
aXcMKYKQSuyCVyG6hfTEx4GZObHNVcs4g0CAHq5DvbYGZl2OdW9jnGaZ44AsMx7eppLlbppMRrbd
4BEhn6lqMA3zts9A3jFpBC6lWNlyMSUze0IFa3jW0rMoMMnNpbuvMFeUHkhljibC4ieSFQEmDZTc
t3WAQuxPRT3HyN+eA9FRrzReaezCZi9bWQo+aTpcQLVEfCtRvUJTkA6J/IstazBytOobTkdVvNuI
o9mt9osNuprUZ3n6tl4xYYujGTq9iQYpFG+g5ISjmxomnL/UJZGxGMio7EulIjCBEfBJZZ37Fscm
MiYaElBychbiSW7Ao2fjQV4qtnsqmrX92mITmoZPp/Yz3+Dql9SNotiartPeqwqsEyDP/o4hTBuT
GmrrOxL4rNFn/UyDuW72vCyic/6x1Fm+/H9pABT2IFCW7U3T/KGWRvlSB5Z8lWBSHiYARYNk7ped
0XZBJMcyAL5YtxDJf7axgYxc8hFE9ivkiD5/ANrUyAu184qZuij2SnIq9mv1ArOTM0d5XsEMZQhz
p/krEahsYtscboX3XFHXXHbAOPUTzmM6IixxpXPtl2ytzgUlEFCyN8dGaNv/4Ktwsglz7r0F0fCo
N7CmIdQqB7HtjXVo/jtQjuhTVjHmetcBynP4vXy/NaPaqWyPsb4/6HVWnNO+zn9Eg8v3MOS3rO5w
JGWCmXcnlncjHBC/4pNTOdUTkJUfFsiswqLZnk2tm69xw/AL69AsZdtkkfP/wIWbk9yF0LPjig36
R7SoOXbGBfpbv+PLKF821DWeGrJUNkB2rcZIXn6+8g6SIzBkT90u49VXFxK/RHa9Erf9QD1/yO/O
odBhboSETRBvAwy8kIjpEUk5ifTh0A9kHii0efLi4p37D73OSJXsMUFI7PvDX5hXDvQ9+kpYW2ol
g/zAZv/SBOomKVSx10yNJHihtrDPLYkF83Qw4XNuV2mG9lVkddrdCpM+iwoWrgHBv9YY/ewWErTV
n5Xh8+PBj874FNEQJcJ1CQkCprTyGTBO7mRWoWha2AgEQLa/cOE3SbRHwK3y7f6Smlkp9gzlXjNJ
YjpwWfGhY5VPkyiKPQtBg8NuO9/MyRCV0irKNcQx3Wm84nIloFnj3SUeD7+6JDpwXv2pBSM4DDFp
r4yNGGExOIaxmb7vr4QEUr4vL4/sn7x8Hsp8suY6IQEy9Lvoc4nKO/462g3Zi8jQ54RcnVTjIlwS
2XEWL6cw54QLDsxH82tTTxNFDcB5BrMqiBOGvNyF+A7YbKzzIJYoCoMWfnYsGftTJEKzE4D/pUnk
cgdseSRe/7vcWkU+fvJ8bgvcLnXeHf2TjHBKADQ/erDOtQqJtYKHijrs3YWde2NUR4Rr/Pa0HroZ
l/nEpgofUYkts+ayAycqFcK/LmNeZJOBCJ3iZPoA9MOmRZZBPoLQ9CO/FENTokjs5HLCjnahLu6X
0OHtnBu30Mcvp0/+FGejbo6Oy6aP0OS2dDzKSumyqo0MHfqeYENZ+4Koe0g1OCIZpbRC/G9DkuaM
HMa5TOP+Seg2WEG3oNOlyvcmOMQiWaqkCKjpCadv6gXq/bJSKh02G7E+n/PL7UvfP4dPglzfzdUQ
SsKRQJHIlOPp5DdEJeUeVnRvZ657Ed0vA5A7rhvGA7RBoIyPpKfFCF99sTAiRGe31kgH4vm0r55F
9dKRSdl4VWQFx3tziWc6Rs4KuYdh5YWGhcBdRN+s7Yz2xJl+ImZunwGcrIb2+eOflPmJo/+KJ3LI
fCl6YjIcwdehvCiTF8R5sw8gUSRmBNhy+hMf1fFctEV6LFekuoKM93iVtGdKRkQv8hH7zXIDwvVi
1zip4w9Jqc6AMwCQeaIb6ywAZamnUL7EJ2qlKbxcUZ0YBm5bdeyW3E81THB0Jou8k/gIMAFxPHqU
p35CCbqWRtQdrL8ZTbwp+uifaeQkMaNBhG+ELTXuDf92HlOUPqpf+hVSVl9Xv51FiC9sillQNSQX
Or+cIt8bFvotTG7gz87IGBgWXu4hM2PI/rMiuwZjwpmBh8sEE728Uy36THUvbt4dmTqSWoN7O71s
fuI+0WWMkeVvJ5PRuhwXWoqj704ydLKzhfgSASBwbwUyJX7Tu7UqsczsCE+9egxU7oGuLn6I6fub
vsN/l8S8A/VceeJHF+BOO9+4TyTZgQ4/VfgezxEXMbZpaYjREyc38Evf43JNS9dFIkwFsXjMUJS0
3nJFI27zW7FeJ8Bhx8F9YLdxvruhd54GhhdGRXe8drM6aDnsrJN8jmV0jWiYGJL7On47Ckmg3u1p
RLNxFoIhG8k/a8LnEyRZ/k6CGeAhkX4FxPYDb1L23z9d7rqWzEp99FqkX5UIfSi6FCF99X+i5QsD
a9WCNmfsldpBMgaIZuq+BPpgCcx/2tAy/xbypc8dPV3q5DeLzGEy2EANsx97BSEiGiNuUGovIaBI
YOVMjdZnqvAZFsARM7gfEOpZvQqQkxFDccusKFlsjecD6qBPmAzhSVfkiZ53w4i8TDoWwaPG+Mib
wak0ov6h+UER7unzwPJnhgM/R6pEuBdoSabaryw78TMkarUgrKjk6sjGbi3pbM6FJ3U5OV+zzUlC
vumHs0rj/SbDHROMT+X5k7yr3ssXLc0TLzV4rZCN28xuW3bzEe17ToUsi7qma4RgFNj9lFToKx8x
Qd6QneXkVl/2c97pku4KfLyhuLGMt+4dI+wNDDN/X38xnq5+BOwijSsdPQmxtjdo21qvglOtJemE
bryIlJR4vJmjCHCUgI88ihybQMItiPO3Gcpe1svmFhNGiDd2TWJ9qXaSzXM13hI8CBxFymuajkgp
fGla+NUwe/8sCP1lMZEn6IxHaAbtn/dEHYMse7DKqlky7KeHm0jxc6V2iVqLOtzaXHx7e0QYaPIk
47JYOsJG2VXGvP0pTeRQu4q4Gpu5dnobciRHlofJlnbaFDdHqguxyboe7EgchUizqXAu3kXOmsrX
wo91rca/kHb3K/MxR0C3lMVU0xK05oihLo+VOrZC/LPNS3XpLwLstrUqK62xVXWkAGDb4YHXKs6S
+8CKPOi+lH9eZL3km/BlKWrjJ1+eZePKcZfE0ccGn+CQX5kycS6WCZI3S0lzIFKYZbAtDna4gwh7
ZzmN/3EWqT4003tqso8lVX6VthH8wnECgGw4dXmin/iyqJ7zjAJ8hpUvdp5nwk1gZE1lexbJGdqn
v2WrUW73dlPXdpo7RAOOsAttOd1I8hnqv089nCR4gDx8pqNMPx8baaI5Nd+Fy5SYI5sml++kjti5
WcI4vwsqpDj5SJ5TvkPM8empbNIqCVNvqa6IDrnNfEr6KTBSeCBrgnZ0AVxOiL0KOUyjj6wkPKtE
xL41EcWv1hR4GHoM5uni6nHNuQCU1fRPOG9/sGdAwRRXj8TE17hHfvRtE+nJDAxZsAxbI5He9ja3
BSNocZJXYnBXAJdB9usM6aaAK83G/l6p+hVkTEUy2F6nXovlgmaf3/ZkL/2GnyWuNySyI3u9tDy5
ENj3hbj42/5dFRR77rtAHBDxfzL0T14q3NFeZK0f8ZS2Hx+cKoGE8tHxP2SVSZkh0yB5tj5VtqEt
ubTMbra89uQX7dM8zQfrbaf4SfBse/9+EGi9f+lGvonwoz3T8bDzfTQqXGPyd4p/qDgl9T7SvRHp
6Uh3niBUYcpS/kwdqHUkYLnQmA3IeMPDuXCDuHq9vq5bXL2klBgoqmUvZ9cvUWmitBN0QdmwCRLT
8PsO9O7S0orEVRzYyB6Ovv4Y5t4qAxx6jo21Cy35y0YggCc+21JJbTq16D5lRYaYJHHFiaCvkmEr
0Khy5/Rnqq/38RcEapAEuOmUkX9VaJXjrSkqa4cEsSGG70vRRUVL03y99DECsQQGBLTbLQpNpxAm
A1Y1Jl9TQH/qw8IceB+IBRS3Y0tJD7roF9ybObz4j+eXisAW0c8HmdEhTM8Y6mbrxvB1mJqntrEM
4L0/yImfLGMF57fY6pU5Ev1DOGLDFOxLSmJprPMun712unLN4zOLvzzbXyKCbLWNtnkQJ20+yGFm
GmCDm1m5SIEqMNGiUpHrg/LVXhlGYTM3Yo/UEVkxiC1dRgSPhDFSurgpibpj3G323W01HyJjvcH8
Iyr+dE97LFaOJJkxb91hofb/ZykCJjymzfEVHZmthYsPcv7zyPUuT96E1lruJIlIcllMoNkRUlFt
0FntJGkAqQLcrpUf1HL7GpdJvNa9zWvZFZ1dnsSDmjnEz9cGw/OPhYAu7I3O8JxNTerv8hFIM9S8
nK9hds0LtNq1bt6FKIOZZLgRNDjYoVjScMnMsTMCsarseKE1GCoBPsLsq5h/9fKxUVn6buHSQJZt
+wxfeZUSyvPNjm+Gka+xEAY/j5mczUxqFThHIbCQrWjQIp8Mq0MIF2FZg80/HDXgNGDxDjcLub1D
gTDuKME4QAWWJf4Q8IBdEM05sgu2t9D21LGJUXRZZYQA+EI1pQC5HylK9EMHth534xQX+hqpbGHc
P3bw+jfvFre+AQMoTRB62au13kepauBPt5vgIx8pkJQe+nARbBivhT3ocXNtYaZzs45xj0FBgCu3
0kSzm/DUQd6X194JyDi2bTnl2XOPb55bQ7eeuZQW0B16tmhNj57kCiIotC2HvC6deTGTXJtnfu3+
Qb/3usiSrL7cMlipebd8eVsw/bSYGxm4ZkIrr8OSZrbFN6lr/GePVp3gmoWH1DBRsedhRjvBeiyU
eK8+gBMFwflhWWKRKyi0LTBj5boz4Qc2hH0+JIbZG9MM1JLSCauRrMUBgATl7y66QPZH/1HKXzha
6Aj8cQ7g5ejeeaVlvttm4HfIDGxAkjadcKJjyOLrsPptliRrKrJGeXemVfsZBGzsaHL836gXuc+F
KZEbP4A1wBhI8W/Q8pqY2KKjbntBCiTgtP1T5ZmbpHY9gRQTStwla0V63F5OWOtNDZLdPK28cwo0
m/iztyxKVf0r+Y5tj4h7ts4j1Kk4TZLOtFVCCi5SZozMmqYZXMlRThYiN/pFRaHKa4uRVGJTNS4o
1vDNWJC85dNio8iGQ/x8ZZCMpq2KcZlvYTrDdSXWfTXPuBXFtdo/Bgvc/L0X3kOJGq7ntbzILS/C
Ngm5fnBMkyxhB8Xhn8dndBeD+y8WlvlOqcy4sN+hyvyR/kC93z25fNxnz1aM+tAY7ji1NFYfc1cA
FVhptf7c9h8TUJydHI85EaHgF+R1zNsN5w4E9okns+2nXuOH951NLR8nXCkifAu37np9loZLadom
jAfwa5DPmp+q0Io9YjMCEaDljvlSu+fZmLXFMa6WFZsXbHo583f9fDb75+wmuhC6dMpwRS7Lvkn2
jM0qdl7lBw4IMmpppOFTioGtxrvrdam0g0Zq1pi8gM/COKvInFwFZ4PT3GZCMZUF6rUDo1EebkoK
EXya8QLT3dC9fjOQJaXxzJk8gj7CRirjJbeBiq2Kyqgr1Fk5WV9ee0gwd6lQ41mVCSe+kIfuqVz3
qXaj+mVoWy0N1a5Ojzn8HuykKGYaDV4f+TDPzY839kNw1HALeHaUn4QubOP7KOru208q76H1zReJ
iEl2mkqfcbS5uTqbj8dtxih/F48zHVpQsoBWQPALuDQzFY0wWmxDS2tm8cLGUJ+fr/u8xT8mw9XW
wackcnslycIDgRb8tlSS5S1f3P4MyeUlYXU9Kqv26V8jKuEzb2d3jVquRvcEoG8ecHRNYp4lapk6
IpdAOKwyAyJZxyVI0s/FX1mWANYAT7e2tQxWkOJZVcO5wJPiwPUCZa+b+MxuF/dgxLzq7XTZfo38
gHp7fpK4enNIDBfzefoDvDu2NafIdghv27LpZTALlFR1IhGbHUSOu2ReJNCq97yhq/gRpor9JeV+
hxxYqSgg7J0vUjpLLRsQjhsVt5co4y1rk9YVafXoTywjnpufwe/oQvTSIfkNDq7yiUutMHtyR646
mmXM0YOQMh4fBqcVecWFRsQYl088eBHDauFBwpFTGslrPYE1JdGe7zCbPccTSWb8omNdLElobkLk
3SvJE54vSC0R672sAan27J0UZON3Bt04hG2SsiP5GJYCL8MjfobYHiIbrfbRIKejqKQPo5JH67JL
X+Q1WajIGnvPkir+09y31IbcMdBKS+KYQwr8MTk9HisasXvUh5Ny/RnvfgrceqpPeXQ3Ej04Elhz
3zRowulTMdtsof0DzSA8LLN+dDp+ctm4eItIDa1VcHGz9Nhtn+XJUxnSdEDjAgICb4HoAci6Hvrg
HXdiFTwe/3kkjX/fqxtM4c74DeOSakVeKZxhWfy1IsdubwqXX79MUx+6rXYsk7+vFHl0FC+GzgTS
2AOaAtvaZh768fFvNIt2a+IFLnnvZvPKbq0Co+PI0dhT4vMveDq8mq00hCmouHd2Q/l4hkJDAuvl
Z6eAPCne/JLV8itWLZaxkSzmcpibAYddcwNLZ8Kf5GouBMfuwXEz+irdd6gXulYlQUl7gtghdjVu
CN4HCU6J6caG95FIQ2R7gia6BA7hxl9jfLhNoOFyfL5smXm/fWVaCcmwyv70tKsmD9gm2vxx0GMx
Cbq1vKjgYrOMTicbAMrwwZbZ/NxazY67VYNl+4OFODZxM1cUrcPUIiHSAFeEpJ2TKKo7uXCVgQRj
pE0NClhxQEGHix/2pBIgPxNkuRkpSnDz11z4k6ylwzWibZ6sMFxnbMGAbM/48F6LcfHzB1s0cb72
nK66Fjz3IztqMI74MNkkiq7HTSTUFUSp7JZAi/qSp11Af4yZocXvRFxoU4oCi8MeW0baawA8QACC
7nNqDoEbAcJ2eZgdVkmbzTBJW9uPP+28DkS39y4Qtb5ZIrV46TWitX5Y/AaODHG9itSuG0PIl6MR
DSjzyVXcY+Ajg27KgER/4V6i08RVqRJNFevtn4BYyWZw8Y/xM0wZqhIDlq2iWxqnsSBNDd8u6WWi
hfJaA28LiuDTQvisIbQsV/g4g7/Wpr7hT8rrpj9rmEooBbZFFBtmz6ulV3exiynSGYeRvZwDvj+P
sxz+daWJLGZhtNg6GtjfEyzoobtZ/lY9qIb9bSRnrOs8/1VBtgD03Z/QhqlYfWAgeD8xKUiUJAby
70Syskoz3oGbZqtl1MOgg/s3mM7sTmNv6RBR27/v5Bt6GHOfS593mSkOQKrcNDdXqoikOXTjtaTg
/XuNlri0DK5SmS1GcyHEcxBfUjb0VjzrLZwr72sjGX3jvH+d8CQZ/aB1ELdUQvwWk7c7OwKvAPOx
XQGlrtYBBt8zcA9tNL13C/Gz9vCQgpxsDLtzQd4hH94KHDHNqWuBq8NGjfETz1HFXMTLpXS8pkUX
TDyjPQpaPS/hDzfokUFk6yiuESB4q9QdfIYYGQdimCqwWZWraLGes0H/0wBe3HxZcoykoHzIM3R/
W+Ckx/wnoZVwWhQHnUK6tmdarA6Jo1ZIFjwvwZ56nI4oCu/PaNdf/G+pz+EDxkXTcDvxCUPvOTyr
9W1yP7/Rar5qXnZVnUzM5W7wEWkYU+uWamB/fzmXn5/3Ltx/Z3yg2vcbIGdEhtCG7dGKdzdxV18r
Bky4pHL48h2SZkUre4OWG49v+gyEmnvNzhPBt12Q6yHDEUkSjSbdp0A1F90S/vZyeoc8YyaOy92e
uJlknw304UNJHwsv/yqVecjVdorhxnhYvEFKkkyDvFlmfD5DUQgys0aRMC1+GqLXoupgTx6Ow5zM
TQjJV8jVWiGsU+6/fIG30ozAgxzH8/FZJHrROBuzSH1pRUB84Dvu94JyLy6YzaArGqZZ7ubTu5mn
9v0vBkYQp5T7BhW29R1HIgyMdrmJaMo9K8ew9w8ZELxgPfTUE68+exgOkhoIVtum5OiwYsCRPC0s
gm9Uyuq9hLyiLoe6xGpJkj+zEhWN57N5SXON+rQLNXaDgK1jen6qhrPFc3wCEi5oM1urgMpygvO4
qUDR2AqiHMLTd+6TrvtGWty4mcchIL5hKzkd2KgOl1Fsr22Pme3Alvoj3WHSF4FWXgtDDVfsVdVs
ui1MeiP0V14XvgKx/nUOFvYlvEnj4HaZd5Ehs24bTvqIwIxmQqUn4V7HNgkeh9j1HWUVnUH3vak2
6dAPvD5yVqS4k6OjsoX9etAO2CeGlojT7Gsp/ylGUNRBr0syLrjQSdGEl914TvvjmJZ3L5xffCKm
0lUgddzE8kiLjf8FxAtcKmJVeX6VTAI20gR7Cxzlclc0Mupiz6hPq8gKQayHg+649cyNIE3Lai1g
GrEh9RRmBIja5vVWlIVptljJwBMwuPRuYCKpq/cot0gzIT7ilrL/Pht96uqN9Hkek40IqB/j76E9
HzFFP8bVQZPJBEUYyhAjMaibt7Io3zD6JpBPmrRRxQIaUWUtRY/YTYycmjd4+uHcgGVxs9AJUHIr
QYVBbNZS5lJvFBCmP0xgHxm2uCDvHjReFIxhy3nX4PyHkxRvTF0tgQlLxkZmbTA/3cV4DtDEAgvd
KpY9PJ82tSbHwpBO5wKhpSBhjTeD17MUJnEPiHdWadP8zR61NRBDE9Qz7VSIokRr8Al4i2dEqvS5
KRTIjraHKzpragZJfnBRGvLw+FPK0ij+/E2aQO/jkWFYUjJKDHzkVbGw5Z8YioLljrpSB4E57xT0
2bPDXglX0jCpSS5NcZ9jXjidBauv0LDkHfePL0HJbWyI8ZF115W3MqkB+lY9XYlSZideqXMIPXuZ
iwotm4ICSv6rhD4E9ZzNNWOPwyV6adr7Omsofb/WeU25T0ybdOJ5GvNQ9RpYIyE4NcMjUQ1mRBXQ
inw9qJIdOHpJRHlBs2GXtn0UtpQabdZvATRiLAiUbvfhnY5dyylQeIWNbNVqdDeaPDV9WJJ4IZaq
PwSN3Bqjer6EYOXZvgEmXYQoCpk79eitbm7W858/rIKHONLN1cHVqzt64x8sFl2fb2utPCxdk0oj
chVmbWM0P96qpsg/vWRfYb+29K26WBZZg7h8lDPuyWDRe98cVuwqIpNktw2BE4IC/L1nGYLweNhh
BURhR8bvWeP1ztcoxyGZSqCVdX5J945IWsirtvhKCrfymxPzFoET/IK7ssWNV6HmIJ565Qw+VaNX
9Wn+IKGG+JeWOiQWnZVnG/bbmaTJXueU5faRmlgM2XxpXPn9lR7s+0VfZoiaAIMBNC4arl6N9tnU
brE/TYtjpCWoOX2YKfLpUmQ0Af/EQ3wV5HBXQEbblwzqzXgGoocDkvu84+vuZJ6ZAVBAoKeWijsL
9JY+ssLNwCZocLsnoPOrI2vKKRseJTrqDmcZN4TDe5kX5KT+34k5qk4/QjvVv+N2CqhczEOCGo4b
wBPnVQAAk4r1Aiwhs/S7ebmp6p+cIRi3vPr1ODGHGqOR9vLqUiZe/KBXsYZYYXb4rO0sTbjvvoG0
IzMCIheorXF8hl+YoN0jFeVSWQXnMLqz430dTl/YdJlLHXbfTONNtlkNKEDYBpi6o6lhsd1AC6m9
m/u1eVoH/1aoM5uQkH65q/zeFxe6I3p/wB/cR00kC0Yxf57aatzdC5CN0k7zDMGWNi6HzmDaGX6B
1ziIfm9amTXXe5ExM/RFomj+JOl0y90MPTn91VfrV6f5oCa1w7spyAM+z1qN9mlbj1D4pVa5+2Zi
PVI6Bvsp31FtBROuozxW8XorePDwHTlJ6FcLqw9XGhPOEyXuc0hODGTWE3P/8EaM9389eq2MO06/
xJEKnqfYfZMdLPpYUyLcOgTMCL48vwbgKGjK0mIPetmCyOvQYyXAU9/YL3U4Z+J5QBt/cwrVKrZv
vqFU1xvPQxSmPqdv/rdzNobgGVuqA+DQJ5mDR4Lavi15qVQS0ZbUEyLjcCe665XxUCSW/eiD0FXM
/W844p0RX+SK5r7ioMvuMpZLiuAK6okz3cdQ4faqXghCfCUBURfVA3Qfzpdy6/vfyFCoACO4sG+L
hYRWQ5kMuZXFbkqpskD7UgSTAKRm8kAnrpjKpK6Ycs3ThOTLpyFy8X2+DhK1dzvjmDPn1lm3pnUX
7YiKiy5eYGtiIIyJqJ4hNi6jeCXRRmlblLDy9AzgOTUSMudxh38tJUCkUbhv2WjSSp3jg5JaoCLi
DXvSVyFSCpgPVeMgTli9M6ygl271uymoqx1Fo2MYdqRWmFjteZeVK2RKJ+1j9PNuEqePB7RW8LaQ
p2hjFBd8UORPNiyUOXpCHSW7uCxGXEeM+9xgd+XDpCROJbl/pqtzT5oG38/aLIdSRle+IsY1TRaP
2/r7cROCvvOGVJe6XEOFM2SUODuWH21ImpDF1eUmr6S44fQ7y0qeW9YnvUNbZr0Jjs6p/5VGmISU
UItKrQp8X7oKSvoB9YU3gsoWNx1tfzRBciWtWU3N4daVsNdC29N8JG7dyaFwu620nlk/KoY9vBQo
w9FAdgI195B0Olr8WzuOyaFJHS6wIzE15rC3pSwnlNuevcYWKOrzvSyqBOkVkMu7qGUONbHItaYX
/Q2R+7/rbpxWYUZdOJnj7LqjhOSNjlEtVjfGfSle6uEeHAlPlNpVDjDgejO/u23Iw/UsjEOxyBa3
bnccuBHXoOfCNda/8H5uGH5ldYfAy7VkFdDNeJVpKpZDr6BM5Fm/Q2KZTPIGprv0I+RMqjPz8CxZ
STLOON7loz/M+8wJ+xervWaeUUhI+vf/0QwBrOGntmevsYKMebXah+5NaLQaIrvduJnYNr2BcEen
4KEz5NSGCNMVOw76798m2T5K0rvTSeXh37W+Yjs/2PAGi/srAFp8xR7GTutxd9ot9+899/VZ2RDO
js4aieyOtfvcxK/uGcD2CTbcse2tiAUWxyt1nlHdwncYp8eH65EZamXPlRqdg/CkJfQAKv7N7uRW
lwzDi0uHXrbM3IZA4QWAHnLKoXvsfd7s7NU/AnDr92zmgnmzbyWTNZ0N/C9zz13M6H8wkF2kXm8m
oGuDmIeacX0UNXRwNJm2Gfqc6FupHr/oCfR0MYlwEQgXyHUMziLJBGM5n/gnO7RRuvkFalfSDoHJ
c2Ff1Tc9PH/9xkpGt8K/MV519EUoJvp54MY7uRgghwbioGJnoxl+TMymh8I0gX2KqRkruT2gx5H4
EG2YzODSCYqBHs4tLHxfMNtrXCUJD4A8pe5YWEQ1wvE9aTl+d5/eiRitP3zg9qihwOPq5oNVtfY6
DVL6GlK/hLEnIKD1CfNlsalb6BUp31jBcITsmyFApNBsChqTwuGD4ZvfLKctoLJxuSaitWV4D5+z
xE4Q4qOrD/3DH8VemN0xDEuixoc2rQFuDoFjcDAzrOCFRXaWgvhdb8a1JUVk0ZgjTI8vdvWrhvOY
AfvDI26znvEYsl77DidfeuaUBqs43qqbavC0oWNim/SEKbh62NCXv3+AB+iFZic30nXjTNpdV/fa
H/5T3vPmBaWnSaosrO4Ciz3dPywnpr4tWF9BuHIZZn9FjKMZBHN1jIP2jKMGH1MS7ZDWQAXDHSoB
+bKgp1wKiLrbjAiiMoOAMVe8M1gWe5x7EYmGefHGO8iJIZjrLL9ywHI/REvqyRnKZnVl7O67KOpV
3TRDp8y4hssm0XEBg93tMV2AjxrfVewaztaNiohTwZcfSuGY9EkWCd0bIcyTpt0J3lIt2gnhQAZN
5NEnprb76Z6mRkl1hXYn0h98nwDfZfi6sMy34TLu3BPV5W9D5lYN4LtVPaL/bXimuHceP1rewLZ+
Zpxl6OjPUhwv+m4u0DnnE08ioIDKXCkHNuk20IOd1gDGOp9ZYKW5HI6JJ353xGxbdSR9a/Jd1x5x
OAu8Pec9u3VLl14OCYyvZFEfDwS1d8aJOmzAoUa6J4rpKkzd2JXG8CuxYlzu+XRitYxyf99SqdrU
IInKmllj1O8zFsw9IMGGLjfpqIGLaZyM6Y/pFXVyrz89etYVmzlplIEqYKHgWCYQLjgJdJXsuTs6
fd5HJYx0L2Q6OZp7g0n48AhvqjR/5Y3GHAKeVpOXUK5serN9OjpPF8/uIGJDUped4MyDuFPRwP/3
mZN9eHdqmDGEg2cmz21JQKH1bBdH9JzkLPFCE/ZooMqOS5QPgR1oxj+ZcwItInBsN3lg5neUfPLB
DsSszZ4uCxqX9mQwGjDZ3E5KS7qiOBL9KODeJLYKdZyNTmjikDjhWHGpXYheNxwhm3925RAduXdZ
ZAUmqsAS2Kn1YwVDPrSBdawEsJB9dNzVJ7Nm9GCXYlYuOXrDj35x3GRF95aBszJzV1nLF4zTrAun
2VPrCj8eTLWNVS+TIsnZEe31gmGdod2R5NZQvj/amGBX9UAOILiFGVV4pghzu2/xaRCdWBtqrDe+
HVjdHg5Ixw8oupNRrVzP/LblA/szCOvmVm6QU1AD8qM0ryKlQfNH1NrySENBHJwy24fwyH28v706
dHf9wgmngUdBhZpaVLP45UNgV+koCUuy/ZbNojgXewFUllWoMeXaN46aX4oVvli3ErrFGFQ0pIpu
q4XNCXQgoW2htvhvsDfhInac/p/9imTY3O2SpPvwdUZJvv410luaeS8tZNXNLoTK9WT3djwDxC+s
9LsadE3bSoWT703NJTRna/aJFSIhPLmDK/ugF1znD2h+N0D3i73yZdVNEDZPqF3DWGuxJHkQDbkd
V2rBYTzpTlIOVmYk7EqV1FDlOZ0reD6voFbu14qEGKhl+eJcrP3NBQU7cjmaJrqPRUBK+cbgFEOu
NO5caVCffTiofSE2qaSCWK8S2U+ocsOr7FsTFt2FHF/wTj3SK9CsQhbJt7xp+kdMymkt0JwGZVFF
O7OqIjzWZ0+RxQ++uFhhhcoFH3tCwted+DI732tI5eOAb5eoF+l2Kko20k4GUryfNXuhk4SwsB2J
iyqJJlhx+TyNArCW2VbWAi0XKnFHFu12P1/GV6vo5SNWB2xVShmlNeEorZt6b0CCTNVHmFE3sWKj
oinNvovWwY103yZAlS9g89ai0cQUlyl85LOdxXR6XYnZsPzMNl7JHdmddMuWIpwWdMYyVTlEJnxx
2pmyQt37HtuV4d45c4uVhxDgJFKgIWz7ZN0BZsqMcCp7FmVV34jdNW3Dw4mcmrBrzIg1g792dUUV
s9zdCqM5xJums6Y64AWaQO0PsrYsCSQebsfvy2jJgTqE4ox24L3hFGVe8SpJMSGLpOiIm8TEwypd
BQh+czQWe++Uyqo/sRc5ZHDoVWQ1E1xFHEKtpLbFZwCSHDTM9q4h8lrE7dyHjHeC/Eg2DeU09s9n
nR4kxYYkTh5B9Ds0tume3Jps9gILHM+Ld0mS6nrltg5+LHLoF7SFKbmyXC8ANetAxTS3POBxHd69
9VrvzctFZk/4CHWl47HDr4zUfavXfmEH23xOi6kX/cT/Q0W/HpXTYSxktOCGu7ddSO0qT9GgGsAo
kNd0Hkcdgw/6zkbRZ3D8hbq2EsKQXOrOB1qFZjN3oDy36NqUvZ9f7rc+myzXrvSBE4WWT6jCFNzs
MygC4m5BKY4/HnUcdW3g4gkZIaH96XovsEpZ2PfGA1ludj0MA6rq3j4M7SlJJQN01h6snLm1YuGK
nM0WwZgHyCr2T5CODHX0axoGTLRoVnldLjrag2iNzJcPBJ9z1ZZQCw58tHeyG+z1cv3OeJoEA+vq
xG+gdMDUiYsWf453uItp2bwQEBCio2Ses71TTe4eyLkU50aB5CV4mbw60xpiITzBXgoVJGoUCBxE
kjrFDMeRyV9PSwP4evPu5pewcLrOzrsAxmuVoLBmXzyJFzp74/7pCknlMxgsv128E274NU1waiRD
1+sN8i2nDmASrNUBSbiab39+vDDaeK5CiIJghjz8flwiSc+X/mgbv98KQIlEZubAY+fCMHSeccSP
cTaWJERghG3e1vw9ByFhRIY0NgX2EQQUVj0y1RCk2BConppHjttsSa0OnzpnzzK6U/WZL9osntCL
VACuCKZOPiIAtF5uXihOiwQlo0Ffi4UMzN2r3p+eylx1sh2TyY5tcsO2MKlXNuKs5htw+ViWnbWn
8dVAaNKARaUR24nBdMNwcQpgqVXKMyHVVlWhMiLz53GxxkXs593X0eiypor1sdRjFb9tCMdmZoWh
D7mBtZHZwYVm7DK/WcFyPZQRQxPetQTThSHfqaRfTJbjtNuXLE+6u/0jKOWR3+OR8gyNysWCtsCT
ROV5pRgsbrkzHZDfA6CPUJ9ccg9DIhu1cwrxbwslKCJdXk9Km66c4iBd6FHMwkT/Yo87N+6pRAgZ
Pek6QufYjoub/4np3U4DtpJoYy94PiH5bGs+SnZbW4cBLbyFCjyLsKuV526hLGRDZiBSqhoFNUdw
S317wOxZjYFwCFOBaE+RecCaJvPyLBNg0NA3ICx83qnNN53ffXMjv3Q3jNIm+L3r+52iOEk88KPk
F1jiUHK3MermrhV6rYLsAiq40eBgZ4AO2zqVOlWflepPRrqCbSidM3BWzbNChhJIEjG3ThGMiNS6
L9a2HLgSWFQII7Ndc1MqGnJaVSyM49XE7P/WXGgxrJt0byLcetDOIk02du65/pNIlxDSCelFsuou
+eLsK8LlDO9Xczp4eHcSrijqDkpppwMbGuSkTMBuVpI5REjIWGfx6S5e87tiVQQWuECZtF7DgbEM
vB7oh/PrhCL+fNzh/aYfjb4dEDB0TW3yf91Z6Ir83qQI2SW/0SiOJ1wJQvy88AZvaCUa4Uns3V/M
We0UH796e3tkCK28pVrtDzGXgnOORPZS1RTpP+tsJCST6MIT+wJihsRNnRgxhIZ09NA0Om/I0dce
VpMYjARu5lfOTJihf/X6oqiiz24ihe6VIKrzfZ4sb47BdZvBtxEX0gasLNXUBm4oHufytJlktHlR
V9fycFMRRNPfPsKNNBSpWo/48qdCWszc7snJhw5KMoGGgxk+W/qYf7TTm2dNuzz9Ci5Iqpc4ymKC
b61OWZXRYTpo0LYBrKew27vqdPMk3xwROqeZBGxBNldIiRtXw4INbtgBDCjJMJZctbvCR+WAOj+Z
HbgT8nLlMhZ3f4o1deD5DD8PeNyBYKGjkxcpmbcTyJ+z943dEFJMkcFKOAqXEmSU4R0NBSVbdgAk
A8KyVT1gXmWAAis3UIFYnfnracSU/XV/dyfhWgWCqynKy86SHBL9OqJ+c2Iq/GkNyP54rt68p3hL
yqRJJODs+kqM1xI+e2y4x1svnhReWXKc9rkqjCGJUgywki0+AsrxvxsO9c74IVgM3rfi5pB/t4l5
+yY5qfHet7+wKBQtx69oHajKMoDgAQG9chv5XObOEnbSgUKTCgQ01F7PUULfRgrK9pyPyQORO6Oi
Ny05Sl03HQ0lw/9hkwmyUsbNGeA5HyECZO0UNV+J8zn2BVs/dqf4uKdZC+kxIyARlNscMIVZLCTF
jrdiPsS7tcc2udfp9WVK7A2pBpnSVFosXn4IfVRXL0twSoG/2cRzj+aP+5IPI7dIdMkjH0Wx1YVC
byEjG9nLxIz//3bZzh495iCTbSA/Yu7HzqvD4yy1VXbNKvHF5no9/nQUa5hwxt/Ky4Ewx0bSHPkb
TLmSeyGkFE0w+iRkePYW2OsWiW1GNcfW5lW5AFwOj+IDUyl2YYfLOllW1du+QrGA3L0sNqDtGUJ5
d0oJ1q+ECM044y7mmF8U+YqxZiyYNZKzFpEHZXrPxervNvKiQRSl6ggvuxZf6RyA6YA3PZFkbb9q
jXaZhlwcUPAcmQUSLj+gtzD0yTfy5rLDgqKKVjZBdR2BIImftiEAi0mvJvhdcl7ffSv/t0BKK3yt
tCUAt/M6mn7si+8+njtYuLoviVc8oKrIZLqiXQIH8gu9QXQJaG+XUAfey4DI4AaNuqcG3adm3KzT
UBv7NqdqJs6nkO4XcCUnMeIMxL7K9s1CRYymQ+Cc+5ydez/sDkpunLkraGe0p0fv161T4VdoDXL0
6HHo6xbkWCbb1DIeXUf8yxttpnbm2cv7JnjWZPzSbzw1gmbdlgrNxyxIgeD0Yfks1V4x/UHJd/Li
xfwvwl0HCbvRuevf5WDEEJiFpQaGLIALY6MLq0nWgoBTGB47kFLduM3zehEKQVc9l091F2VvEP1K
dxp3z0vG7JpR+4ohb6rkIar+GGA89vIwcmMC83bylQsUdPz6wsZ8WwUUtqoSMNGeKtykpSTN+Ure
WwZ4nOvsEOztWMhezADV2pMYyVZcmDZrBv9MQQDx7Tar9x39N/C+4uLrOLGXs+XKgMy0jS73OUcd
FT1cUOcOI0jHOVWSvMo9T0XKcrH6OoUAzIiuIXxzTtGwGeVPFA7BEsk9IolTgvO2hApG414tLK9Y
+8MBwL63Qt+ZAo75HSG2E8bNt7zmgFLDIKLBg8Woj+5u6GL/hDpOmdugwvZobQPclZqNmDvbmuuS
8raUXZgyRVxa+MEFLfX59Hbkc6hBmPxKmcYBLMt3zz85u760VYW/Fk1BYGLePAyEun1YR9KXy048
B3V4MbMRll6AcRJQQ2ElQCL0g4ZML3XBUsNiijNtY3tjPyxx6vepWo+aC08IADTQD0BETn9DlqqI
dSb26tbf66qP60fAXU01iTrqIMr+uleXyz3uZtOywyDi8HtdW32Y8Z+0V53D3cbbbdhEV0DQdLCd
zCmmHDg+Htq9QFF4NUey43e3ZdDm4SnGdh41gfyCpV0UDTzQcpVijeV7rP5b9NyBRxYMVQeWymhX
KjkI88oBMQZH87lXbmev+ElFRR2HWm2FgCscrDVvg2u9G2FR7o3nl3wZsV1MOUcjGsn7BybDuwAf
9rLyqxC5EyCyd8MVpXQ+lVC0Sd5USGUZNbnSK9/UEVE2VvKI88rsU1yXtv7ebsoXdYB9jDKncPOR
7hVoLkJA49+sl0icBkFnjDSFRwNjb/7gjfWf5qrjPZs8QBcON1TvxXmDZKDWQs5pvSzbQ2blzgDi
F/0yacHW8okP9Nn2jdVjWPlUd+tkIkuE4pkOYRzKdRTAwIJhh2srM1QUUcCLXTfR3x+7Gg/saZD+
q0tQ8Fd2TZVUhCsXM8MP47aM5h22mnZOrG9Sir/OPp8qNE6Lm2eaECHsJ0uOkZBEcOEM6456Ha5A
EMwyfabnFwjrVGHF6/zOdJbTn9HE+QnwwB+eVZqiuvNE1z+94T45zVEHU0ObbVeKSUAfNGn2KdfZ
hwUznSmqlmaJcgYlwErEQMFisSwqINomRsU8ELBEvBp/uRE0GXW3gVgsGWkTWWr12CIzdaxGycXi
4bqStgvWaS3Fb1QzHFuSd1T3CVQkfEiSVMWB4P5+zfiN67KKHSQ/T4MuN70WwQAFPR1S/rPWbnrU
686J9Zbab/gYXGn6Q5beIj2oAgI1kfcQAEO9lA9/uzL4qNcbHuiGQuGzxG/6Lw3A943CdGyAx2mM
RUcKFSSExo6b/jJ7MkMEC1YTgVvlFDT/4E1LXfDN1VH09hi9mWCxCvUVC8v7KFF73LmhNv+R1qKZ
HOHbokFxBu1/YuWg949c32xQ1RR41El9pUAkDXOMyme4v8ynjZE5hXdcEs9u2wpt2kEvTfHfOtk/
w/WMFtd3VhmcZg9mL4rS28rdFdhiViL3bqeoERyBEwUPcX1RdUYfah+8YS7gPYcz74ltGBrDKsiv
CEOblydl6aVINSRVOkTaE7qev9tiBz3rRdKRL1WVWIGbhlc2aFyZh5BpIc6VBluSuQ5QtJ2tliyV
8jpgnNkP//XXzxLpzHGlGxBq3vXtIt32aXFaAw8/5+j3N6nYIjNcOa/goR3bSfwkDpza/OZq9cpv
xT8zussjtKqkoMrp2qn7ARb20ifsPve8a6brs1/2eavmYpc1w3JCRNozE/DecmkVO6TENaT1lwY7
tNmo0oRcTF+QpKqKnS46axQlbg+FUh+0BaQI1YV1sP4TQ4k09LEGhmGoQyZb1V5NCZwWRU2kY+9q
0kUInGBc60BeNO7b1y/ZNe/PgnXFA31lTp8KIG3MCeRQo8YDFNnUbq7aM4Fwo6G+G1bDMLBv5TtU
zInZL8E9MimpIOMF3gNkEGZkF70PMtlPYlMKnEHasPJdlL8uYW5+W9gQcXeA25GTihNFLERHFv4s
CoNrXPu2dapqdheHMEj5EaBPGQlxqJTfgOu1l3cx1UBz8wIaLy9hbwhuSEAw9A8weZZnRbTd58YH
+GiJbh813iCxWwo/onWKNzPee4xe7qmJJ6r6BOHvScfad5gH3iRd2SeleIaA/BWpa4tSRuDX3CY4
m/4tgPZ5Wf2Uw0igBR/OBtCXAYU7kotDcRquAr/aQnjF7YvziUN1BPy/rAHy2OaBv/AtFs2CNpQb
1UBexAiH7nQFWD+OHPzWXEFqDFDZIVllhivkqZMcgLTeA7Adn+lUyYwbPgmjyxq9+CmTJy/WaK1s
GN6rZrKVS/DS+1328P+fou4/t8xga5xANfts6GDMnuIIjd+N1DCGd36KYTV5XTngP+bLdIyYJouL
rrISUgopf3ba+svr7qagbuAnG1lE9uo/1/2IEpwTwnRWeP1/q08Q/Lm5hu6m9uH45Occe1VFEDTl
ypq7CIpcL/r0NjYxbs530Yrwc8StzcNt+Lu1GzXDXwRzCyibyFnWCxr9gDHgWASYAaQJAF/FdoJg
nhtAk+ZUDyFfZtzJlt/DZKdG89B56mUcxqIPy+OIStWI3vKU6eJ9jWoceV8ODfuQfBrG2GfrTtfE
c8K2nTZ9vikK1ao2t6ASySqKpDXQtzI4T2ZxKfY9C8v8v2Bcl4wAoC04KWC9ZJd9vA4NvMd+7RRN
Xa3g1j7SaHv6sdW+QN33Mm8g6JEvgPo3mhwgyjnMcBsJBuT3OrC1LLmbHNKMDTfz0eSDxC5opAY6
EzHoWfZyMkoEK09jKTbH7Z/v6f/EARuTpu/if3ZwssQTpwOmaNVvmsHnTlOSY3lID5XL7ur9Kj4h
JNmre76RssweFdPcywRRxqv6wfYjqJtAG9jNAXKhorJ6eWGAVLFbxUiNhU3YISgX/RrUhhhkxJM3
aAU0ULcXpQAefXHFdld97FN0E6rySL2jEwmhcVcTy7YO4jONl4Html4snIUm2TOcRh0ZInJwO1pr
Mr5AmYwQ3M2fMNbAbCipzmWfvFerWaBRg0MtaTMTdV/2NR9OqdpGx/pzDKOeh8OzfKj44IarYMVY
hMdUErh8A9dJldnPqHgoHagWsvjYvnxD6dHlEM231fgDQiraMT37wVOJNEzPPaR7xpI+dNR1lMaD
djwAxJwLLWGlI9HyjdAVTMPkp30brSfBxUhzlj3Zt4gNUPpIsxDbR1KjkxqhLuvKu3yQRWp+FFeW
FIuyjnRG2YN65KyOH92GZO0i1jzkexDo74qwfufdCOuAorWwOY9l8+1kT5a8kY7cwBk+CFnwSiM6
RB8ZZXI28LCOV/+G4ulHxhsznxR5V3lHPblgxHORm4vMzbOd5gzL1KIt7SxuyFze8tLH3t4K4e1b
hR1MCqHYZh5rS/teYfzk+6R4egO3SE1f/YQb3PeasWkdZP6P9rFuEWKv+1/rQVeaXN1xi6OJHtNv
8ZnlC9ZGV8IB9f4zbHnkXFW9FLvjKqyLSck8blSPL44IlTX3R3FutoOsoxQszl+YbT5vIWa0Kh5F
UPfKiKwhWYdtrV28F4RXDgFYvBdarqQBrqDbBA74O4KnIfr1Nf/Pdt+5ciWTUvKbBfQwtp8l71qq
kO/1Rl+QL/PxkyU5cDw7eidkmFLWYbx2j+QChcwfI6uQt0e2WcXMBiqpqAzDUfs8stVRTSOUviLx
2CZtMnAp4GdbcKfX83LWHReBfv7TqT7G+2iKCnn1TUxLE/cUu2cl2PSUezEtO5Bi5IMN224jlf7k
ugC6aIJdqJg9PPoQLEaSx+OZY8HX52FxoIMWVcyswnLxLFcrYK6L7zBDgTl2LDoP95K8kSzpzQY3
XbSJYELRX029DVSQmceC3dL1sTuK49N75Th1vGfhWwX6omehZTlrxnOAOhLtARuQL+XGrtHLHFIa
2KR5mbBo4Ubm8h7oXae8jYVQnQ4JPfswY0SCUR2q9J2PWcH8WENWsXNEL04Tu24qPqYdam2lQbAK
C0snc5qfNZUps2Jf6y53EpNzefc+Sau5csKeij5T7e0IAd44APoT0tmn1Unb5kKIe9CIhFA4Hd9E
se4wkZKpj4wuNJY7suyiPLonI4WrhJVXmQB49yHOoq9nvNqUTmWKjZe8YUu/c6B8PPBjvtJFVJ66
TqrIXoZ+/AIZOydkSlUpR1wz7I/eQUGohmaH80cUooqsUb4YmJLDUq7/o3igC2BQiOaW0IkTbsnP
l3rSiGVk1gf7DBofScf7DmhQgJ2J2O9jgZ3UIARm1SRuBVo8BY4FS3J4GGnQhtmnOJAJRtdFT5tS
QxXXmYQmjNh65VaJ80wT9I/lSyVLaTskDA1xvkLX0zAv4iewhlebAgmwLbTgarPJ4lqhrhFrK7k2
sSQLw03UShLxAn6RBvKWyYQ/+K9xuLoFcQ64YxdbL47sltmsKMfjdp7aXIeRZLiiuIQG9hl+D48U
7MnFaLd06V8VIPdqwZFmGANpv8Ihl5wZliEMvPNJpz8ZhYGZPO8ws1euaFcXjwoC9NS1EdTya9XT
Q+OA6dzwXXfeAdgCkxye+wOAD41x31PPuivWf28Xd64ovvsA4j6Zw3MsCNFNRHROEKFuyyy7ADGc
o214jnwNy0y6jiiWFomPSTC67WOXX8NBV/WJCM/PIBnhcS53yaqy/C9YlfIflkc6y5JQH2qj1hGy
islDn8bnZ90IDX5l1XCF26RYjfIuS6GLtOIbo4SYfCEtgH3WC+jpxefPDL94FhYAJTQmkjTfVfJE
Aw8Fxeb/Me23xiU23DYvdTFpGaG4b2HKWOrLYOLcGG8E6RkQebhC7wKBa9TfILzKMX+ICbmwLV42
s1Vu+WM4Ob8lVuQ59btTjf++btlsxz84sPEkC8CSz/lmGngv6NjhPfNHb/A7ZWG4f1N0z442aGq7
9FW8BHg1RyuqvXDXKQdTwGqx6vRUkytzSBlfUKDs+qWIv3cRkddDCmbstveBpyeJoAV0piu8C0Yx
FKxkxtGOMq2AvjpZsV9CHrc68VM6D038sPGJHwdQb0R4zaL5NIfEmVSXy6N4NXgkg003znT6HtZm
MeviQUm7jQSWFuntd+JbkzhTiceXCcrMFV4ZH0z6j5KJiSqjTtwGocfeEikmvuwfBWFBryVmv1qc
OeQUyLMTl3Cb5SUet0x2pdDc6ITvg3uL2KP5tyX8c+v9l4HXU68QdVIQbLmumOwkbLj1YPY1ljsG
6vXk5kxbAAxaNARUAixUSvkJ8OU3dlmfb5DHDPekfeZe3Ov1s0lCBT5G0ps+tPENKySdzKQFQePk
781mpd3qGkvDozAFOw46OuLuif0IJu8oAOrnKOJygomMHxxoj3Oqlsl8QBzS83d7Hkk3FVVMcbhu
k1ldRHokKKrte0iuOpF0wMdi0D7aEd2rsJALltBduNReQc2aDgkyYLpD7Hugs80XKd8Ntw9hHr5a
uTpB3agIxTsofo/MNdz85OTDJ/nsp92udPBY1P1uudZUYtPoCIbvzSj9P34sjD/Sho3mrQshUvta
VZHfDwnzEsc32OZIwnbNptvVGb0h2xeSjvAojOutxtc1oV770HTfkANfcWGls/NXCkv0w7c/NcKP
nEi755VrcXiliFIMMGiagHqd1ei7fzARU00hsUV1sGkLGROyRc56W0gkVGdkGuWsPgbmQfjGrOJJ
byPuxdag10dfdWO79R9DFFltywbq5/fHgHAl+MnjPQx7KhHPIxnJF8UnP2KasYBe8D7EXDcIXIDE
QP3QFr3/+kl/xpeQKkHi9bkkWsgkxQ2Cpe1+NmHnU+AaN+KUCqqGpNXbGnR9frQhLltWopMgHGsI
TDub6Ca1zbvXNy+NhAHPBsKL91UlmcWBDZQDyF9NlXte8O51Lqkp9j64y762Gjo7yd35B4py58xY
Q414wGbxlz8heFRUkR+Cs3Ka3dfRvb5VX4RBhx51Nb4+ln5PNDte1XEa3wgJ3hZgWT7RrbvUP7n6
2DIrXoWzg9nOznSZZzeXjoRG6L8/fHJyz33zhA4mWzi3HLDyXZcYTI1PxG2udmCGCIha2rkOrB/8
ZUpIiI+RZQUUUnFFk6ZUBZP3nJTlWT8n922vhNvEdb32pJlLtmoXZnOXJzSIQZYzz/Hs69G27N+0
oo2OjmnGGSL2CilOHYGTqNJY4KCb1X8eiMMwGQ72nzRZ9F6GAQ+JImpZZZyQxosw8T1p22m3SiMj
aTU+BsMOfqxxf+lUVcsNnbvfIGjO4bneqSVkuWP8sHM0Y7zvBdFrYYokoix1dI+aisBT9mQAOm9O
l7jHzSoGarUVW2Z6+7UkDc+DTcb5ssgIcXG9yJtP/Adtmew6ughWgETIXTbkCKLpgKp71hrTAYg2
wxrEcABkXCeWGiRQTvCp/xcKdsoNbVyW4ByOnIMhXIYL1iLvCQuRTwbkNu46u/umhIXB94LLS5LE
AdNu9v6IysmXAgZKmP2m0/hph5bcVZhPl/WqKZRB8PxwHAAP101MFc9CzwbHW9aLsDdxGpCEAt7Q
14oQgYeOJUB+jnaYcwPH2bPXtpz+i0M+n0QVyIPpkwIGvciWmtj74wFUJW5z3IzRw7Fl3OINImFT
klSH2LlHju8IxiTl9Ws6MEnxjClgWRg97Fd23tO612MMH9TW3vLmO6XXi57fTDw6xPMtUtY1hOmV
l3zGskMDeZAU09MH6Ha3F2xSX/WrYXAfjyvb9HuzOmaeH5T5WSZJpJI7eqt2WFDosXlZ3zRfK8LP
lubkmJ69c/7uIDG9zxi10w+RNxYAZy/VJDgwOOfLPJukjTNaaK6NU3F0/H27JnuEYfzmn6AZdDDk
yZWQyzKrgOkV0L3P+BDdGaALWvkQo1Q/IhPS3695ujT6OA35TZLGpcA9G0i6Ee+gyz9CLBqb5ppC
Aon2x4gdM9QVE+wDX/q8K8pTYUnIDYcaB4e76n69M5/5mfyNBeQ4Jqiajn7KekKdyDRORE+/Iv4e
XGyRpC81dYX9ftlEAa4TaG5MgUTieQtDB4sUjR2038+abndiSGwrsnuM7g0xe64pkvF+1BX9vO1c
5Hj1p7ElsLFr5rgQay6QMvBmyYgsNKXRh7g+/f4aIvePoODLaoTKJq04MAcG8SdpxdHvP8V5imN8
BgDmRYiylS5gpadBWEoGp3gV6Dic0Yqv+7Gf2tjQLRFKrWSevV5HXUraHcL4ASKvEX9vPOUZCdBw
odDg0o3damZQvuDvBtKvwKlmKvULR/vodBGSpcL590/XTPXsMMJovEWG/zLZ6IXSPM5Td9PrD/40
aM55GAZ5U1lqUJsuzxHZw+lQRNggQahyp2HiReK0fL91+e5o8ZvbPpniS6po+ZzxmOuPSSAvMJKw
5AI91XHsdjiv83/6EBX+GOfVLQ3voLgJ7+szKdCJeGj8y1K5SiF38ra1X/PvxMy8pMRiMPf8xj7n
V8WJZrIkQyRAWYbJbfN2Y9sWr/ddYf4bq32qTRPpKn8sa/oZCFe/ppf3DfZupTYogFuH07ZAJ8QV
HwhmbDVRnhcqOy7rBQ/V0D458NcqK+ZNTRp04qUHs4KiyGIYIwMh+pkJB5SxXXofGCZyREuZayhu
EJtLG2ibDMReXwOFWmzAsF8CcN0y9Y+UTllGlsfsBG8B3vunyZCgnFVxomxCucY/64KDrQwlIDhy
evY4D4CAFVReLmIwY6jL1HOqIrKByG9WQggC4pecVk6oMJpcOHQ+lQbJPNYdxwSsfJYBDce6pP8j
LeBFisPN7fMWBJOv5Aqwb+hvKmuJR0GgaQAUxai0C9eVX5CmAc/aBaxSexlQwavho82Y+Oud//Lv
qZNFicBO7W+padUdTe9HTwagI9dtA4VR4iyczzWYCElONDWWEvqK8iEyU4dWuEY/UGLzPcaDLiEI
XtPVk6E9RgnQ0t4FoKdzlMK3pGtR8WLZOCPxbt7U9r/jAmnUNFaM9mposDX/BbpX1DU90dPRhU7K
tBMSZo9Hwvn2aBqIIVHDJ5TXcky2qKKF6Vrc/u55m6GDtjS1cBPvtMi56/tAbsRtmvE1fV62sA34
kEE354AEzp3ojFNvI24cjiLwQbsfL0v5Pe13PYvMK/J4nlzT1nVt3HKv/qaIwXagAqzLZR/rDafy
fCeGgfO3Ap9MhSaNIXZdiQ/JDr4tEnj2GSZP3n7vviiog9DRwls+Yh5V3Y5276bd1LX1NtsYahVr
w6WUupocSO1cGz343eY2sAcAwfMRx8b9on6UgmUK3RoSzKxaN63AshMIvz/f4/GUkfOX4w744gi0
LVkR6bFhLNQivMAS67o0CXRRq2o9y0a79XQvulRtE1Srm4MGlKD3/uvLsR9zuk++/H6njygUhfSV
AJeLH4EXZVAd2bRw2vMN+jf3Gx3LNmAfG5QdpE34mwiVxspSwa0ZD+KF9RM3Dz9Bd+pP/U4K4Og8
boZVBPlb8a02cBxUeaJIWu5vL2p44Q5UfZyIOTdKddJ+GfS+MCXhIilsMz8K7D4lAXUMXxEijboj
a7VJhdN+rtk+aDOI2OlJf3JE7CwI9V1juWEIxUR1kuo6zzXSEvbLPEciKLIYHdZ7QpussLGyPevv
g6pahlgq3qquvWWtaaBtBxcyZeYZFx4bIKrqRZaawPBQSQBdkwDGOApKYa+IzyxUaGwswHeqVgYN
Hfo8KK0n1VW3dnqdMOMg9HA+r8U3vo842TgcUG1CuP8u1DDapXFNILruE9xxVaTQ2u5vaM7vstQ7
GXDoLe7wtSUUviTibQG80wQ/EbpFRw4drRAoxCk7JMC25DgTLQQjwhzclh6XgNtnhyUGarJ7x6I6
DH0fhfzYhO5v6XzlpoQMS5aLo8LMY6L63TMAQbFNIsQ8qPLXtH4oWJNjySSozShVKuVipSDGI3xW
8qbUT01s+dl1GoNZXpsT978qa827Jr+hSGTiR0Wr1hfuOYdvZiyLwuRMVxQTJJ/qc3Zl9ip9+y8y
+qA9qqgh7f4gZTeDcIsT/OuXiSLoFsk2UryHmH5DL6BmpSwhiyrejFBxErEDAeR7mPC0ADRrS2lS
zuUI0koTcCKPdJsGpdIJaih0lg4JOhvYzT3b+fIlbS6vJU7YfaC/0Qy9GzMdghmKmYZ1v4Z0rpm2
sh8fgNUOhAEirPv/HmbnnzKCPZYQvwiE6nfOscXB4kTWfKhp/5Cs7jyQ47tJ2fjokM83P6xQXFQb
kjfdSKw7aQTIq9K2Sq0aZ4DCRZsc1WhFE/9m7O+IAX0OzzDwODvsjdLsuTe+3d9KI4epLLEMABqC
CCZ3KxVQbp96OxX71Qysos1vn1KvQxxR3EKwbSnvp8iUDSE9l9UBRYIzgwVBzym2mBuBiqTlUGrv
3Nq0Fbskqcii7weqz4yYMeHlzGnqAKJEiJkE9siDoCYy9teUox2wGDFyttJ5XF6lx81zCMrXSWEo
9Bjz/JW1lUeAKKwF2bNeNaSsw6JV61hX1WqgbLX6a/ikdsdMKlPjH9ZjLwys3LTWzs/7pr7vk97t
T9ni/d7FG2wnm5l6YnRi0pLdZZoIlwzoV0STUkV1iQSLeddpXRje3kpwH72qXxljfQdbajXUNbVd
bhR6KMRwga77dP6x9BqEcyLbzpKLjf2g3hu9xd3HOLOdH94dxbTs14cXkxbrcHKavOBVzxoT1/+c
vKpsTJmT1W8x8IYFhL+k98cMc2Axxjc4EbVJT+P/7MYw7l2ToUsKxmxmrD2uMMFTHuBaNqeHkV5h
R2lQ81zXFRPhQMcdkq1/5maJen/nl0IIjKv6CRyvInedyWJYjli6dfnNTV9fh/mN9kAKyM8fHmx4
pEm0MgJI1Ed2KwD0qt19UjLlpG3adDTnREz6sYkuDrv3qf+h1FwwuL0JcbZWk9GekYfGqQpAWOu2
8VQjnBLu5G1EuS8cLhrYZGl8YD08xrmLoWtui8bOyz0+iwFWJBhoOAdw/F2xD7FEjuunxIIU4mbo
C5HzSVj932Ghehng8h2bQWKicx+h5BUwPo18ZkErncGyQYUQvHrP4eP1QU+79DL4l/5Qre1tkj32
yx38neeRsher3R+C8k6JK4WZ4k4Unz07mxamFhTPduobUb5ORuS9DWUPK7sTgpL3Mdam08HMwr5a
8LK5AmUzA7VUDWnu+Nqvsg/06V1ZsLFF7jAEoPaDgvBR6OumqGkV9zmQF8tUTqRrn8DzzX5Q8a9U
cW9EjNw5RTE1uXrMeWND6BDTHFGSSn3WBcHYE5IKm+CXCg920NAzVVKbl1Yo651fOCvivpeg5UwA
nS+SsGzoQQnzo08JoHi2iHsqVY1sPUpoOFwXPMLMjI3u5RnONwW+JJb8uaniqayW52+X2tjmBeee
+rI0T1/SegxTR4X/CT6bTTeGGfLCDbUm9JPujgli6obWtOhSl2p5oCfdR3OEbLLH7bt7ZuRUqYFI
glicOt6QLzKJWaJyfkSpRa6S8bE1oCHTFsbxpPRbVgfuvMdw2WS69f+wiAnBjkT39dS/8IOwTLDZ
Oc3IB1EMun4w7Sdrs1775XRG0VC+93xEmSZPqUDPYRPYw5/Qgzb09D5Gh6PsXeC32SXLCMg7/L98
gUGcYAOa2lZT3XgZcnMuRm41lFudIui9gyMc36m6xe2pIHirGMdVdUkbu0hEN3AbraZrqCNYkjTH
2OLVQDwlSSpYudWWqlYUEy+uOdFT7lWuZoAGRHKoVG+18zE/Ns+YyhMQ1wDST0v3OLzutklsLsdw
1e9plrE1JdjU7eLzE5p51WAvB7C5TTdcm38MDHZdVMui11y6F8pIDcjSSMBDvXIAqZWfZxua/zd1
1NY5CvL285aULQNjsQnTRAoV6+EX/Np8YU5g6ade8VqPLfzPdfuHea9kDH9LBxexzcM9jqpuxU/0
UKr73HgjR8x6nJBsI4Z8CvQq/90bAvSEM5M6rL9T5bY9FN9of0zxOgfr1DT+o19orO3K1Pkka00E
FLPrBv0gllrrvJNyXqbpfbzeqqU5m97Us1QD0lUiKCNLMw0YSbDbHM6RwaoiVOhA8hALXQdeJQ9q
hlIEikr+hE8rdlKFOIVYCr0uDwm0VldyHFAvMSkLBfSTJlKWFGzFvVm/ap63FKSBvbypMQLhdRuR
tI2KipIhMYO9u6tTpVsJgYqglfPg3SIHQRjQX2Jk9ATxQe5s2zL+adOs6C1ijYr0Kr4v2N4ox7+G
BIYs8crAyfbcZ3gww7JV6Zs0FaIw2rxOIKKXM9/Xva9QTLTHmm3iAdrT+XZ0bDv/o8sBk8TtJ5J2
LzDzz+yhGODEojMck9PZO0jmrDpbWPBXLQ1cs49F4k6bQVxTCQbfRuAzuEbpKcG7AU1kETHpTNxW
yeQLBJusLOcn3hz7L3S3J4cvl7MBli8nLVPDPfHkX6wQ5uLZDUNjxlUL4kq6roEmMkdYZZVCdTds
dxlAdDFTiOi9oEs8FKQA07hdrZXs+IydKo/OD0+dsNtKK6DR7OGoiZa1ShrqVwyg60DczigOENd1
AcT0nnRYBiEj1NCMl/K+uixghAQlmaFqjmTsq6GsDCvgQWQxf/IKcoUtGeQBzjv2SLEKDlIO5AdT
Y0tzqVU/MEEEQarVffPc6976koNTO4HQnYDIsehPKYKHyywOdt89Vh8I+/QHmZBAXCXrJk4C2+GX
CgBFvg2akPFJmtp8rbrN2PyhhGN6eM5qQDddikPrvzmRV1Vwt1bRVLTVHnQpc3JMgY0o49Yl4MkW
A+l9zVhi4QpYJ8o9YuSfIpZrDsJgZOGkukElBjsOjvm6FN/17teqWS1H23S7atvmkI3btsHEXaW1
e7+wQFE0p+YoO/ZIcHsJ4yW6ZjGxjc54hoD+KpFE3+Ygx0E3fdY4YpxoCR/CHbdSKodDIs+Bdk7q
AnVFjrkFi6TfklQpREmJi/P66vMKHKZyfCr8YkEV87UwISg0pwKiaNKd93nkKtiopb4OyaEnJ8nB
mlFcEvqIuSgezMdhZWuMI7pnfu+opxnB/dvmtlmSwvCXBnmd6pnGWwj33YBgs/MXq9sqgInjsaCU
9RSpJ++x7ZBw9txtDq2zkOcTaAlsTHaL/Y4Bl/l12HLIhobb59eS/EDb8mxFk/AkmUUvp7cXlbpf
b0VCF6M6Qud2DUXi8GZn2yP98NI5mR1R1aumtiINdJNDjjKgFll8sGkXyLeMb57xpcMcNmRmdYhS
6H69xSS71n9FH6nkXGmAp7VojgLRIxy1ZyM5JNUHR2/ftqsUhGbT05L89KyTMNIkUZ6nBohvn9xI
xBC5UsUNblaj5/FjzenUFB1+X+j3vCHTdZuv18WXc2+aQhRYyCJkRu7ue8sXi6w2wAyQF9m9whID
WtRd+1a4LGm+7SWEouW0a6R34KfVwqtFrTYA7LcW4r3l1zvKHUCmo6PVQJ0ZHKNlZvQxwufqylh1
S0I3yt9G/lcYLiM9uexYRT0Zh+PjtLaDc1BgUvt6SCz2wi8aLsMLk9cmlnX7NKntloA+Y7qEckkg
+GIM5Ag50QImS19+NA1ol57BzCuTSLL6vK1nEG2hHpmvJK1rKQHEtFKqmpzN0HHFaWbvyvfe6uSi
1L2AlJyEvfozqbofpgkkwy+XhkoVPtL+wyqRKA22FS66ogVTjEYT79Ut4uhVI/fNajrwz2o/Pevd
ov407OxTBJ2/JnpCvVhpV+54820ggp8nAdlIdPoRaYzzTK23g+b/OKMiyVDQQCfcMQ5kx+YTO5BI
TZV0u1Mn/2XbrLuI9SbPoYpYFBfsY9Umh5jPtWWStN4DOEh6WjT28mpitydJDHElOlF0dNHMsGGP
WAW3nonFpIlAYbG/8IzwgyGdcSRZ/X6Elz375G17vm708ehf9RI6MRQd0ZQIpVp24wKA6lJ/VYCH
WbkZPIN46S1Evs6VfIm0DR8oq72nxt/1m6v8iqlgqm+aW2iRc9E5Q7O7pEPhL38qk9IJfA3s8LIZ
nDsO9qFykXoNPN+rY95CD/w2/9IHhsd8fOlvdDXsy7BZzul38as2D2OiFq2g1JyBVG7A7wTYXQQB
nIhLmDEvcgh41nYkymrK3u3jyQ9zxSqtkiN6oj5N3jp8uYOIJQtwvuMk1J+jdxfMk1VaDRC66zgG
7/Z0deLZNf+0VuICM1aE2W0zQk5UqJyVTBnrY9gz6KE4DMeFQIX2NMYZKSfJrFwxdjjz/eEXPbjg
e683RgkS7+oyHq0Ppym9DE8nLJlJdsOn5hUggJLVQYY+JLF5NIafkNjVO29DIIM7mknpOqYbKLuB
0MUahW6IT/BRiBerBdDv52xvyBKqcWaMR0F00SrD0HUYTU6cjWLdVJhYCXi52I6Iax2OUGD1gyUR
CESLbsIFN0snu8+f2AUqqLVGeEHWAcz9slG5jw57ijKC7pUqKc2BcQDedRz6KRCjmXw09FfZh3/O
uWeac8kwrPcmIh3b82t45qkg+MJYfHI6yOHK3qPCH1ty1Mb4915Hn7I+ZpX4WZjwAvJNzDRtWj/v
d87A8KVlq9JPihDDttEaTkUKGO8k+qXF/s5jp49ol1sn7emMnZ0OsX9O1VdyKLHRyyOytWnMzoqg
h4LUeD0mEsbOyl0XeQXYReH171clEQaO+lzZmidcIbfvqBaIYpTQ9OvTFLN+oUWZ4Jk/ewx73cnG
99UY04v60mKS3yScYL8E8d9f/h3tun0DJnvH0nQqLNfKPPQXIHaonj+6q+bg5qKjcXc29MBYYaKF
0+lBj2rJ3L4IPP4/0xhCAKC0bbz8ehkOQzmmOunnj4xnNPjq495xsvsokCnrxXJiTtbVN5lb6Vrv
En70XqstjIY29v67PjQttcPZoqcIG+tGwg8g/6vJmPU96cu1KCPh/V9Wbcuwa6o+5VPdW+lIR7sZ
vQItG0Ckn+Bqjescf/gcHqzTlh8p6v5lWB0IK9w8wlOOcaW33FadD//wxjVyvfGSKZekLRQ2tJmn
qvRMT9dItcmMITE5F5kIgB/ocokQTGQAwgneahXdEU7wYXTmpldeqUxMVWNmjgAhVlzzC+T04N9o
ksMue0xu3reeE00+UH3UQDcFNWIYfRF3wRouPM4VZ81ddfndNOBNP1mvEJdtPDCBHekCw5QLkA/N
PzaOZoTY/jd62BBTZRUccPfnOomdZWJ3kpcTIWqTJam2jyOX39Tr13RBdVw/+6RJkcg3CG7EzdkP
qRbE0EZDHLEaBgd0MGSYuonKiyCwi7niobog+iQui6zsrzFZEYbaYDwZkB4VajhXKHxIUjSmEcwd
HhYqd+lqLyRoWD18u2Y0VN+z/yfXJDew9yAn/s2rD+6rullZuz2PuJLzTyM+QvooSQA2GlZCVjH1
HWdhEw0DVKQP8ZQA5vV2nZ6U8otECro2MPZ6XnjMGEjosw5Uc5CZqiA9dPCzFFbFCpGN64NBLcFd
wfpOS/xRoz2PXGmhipoXLNyNopu5zhUFHwNxZQpFlchjjuR+n9elfFYHm2KYdwkVNu5VnIEyxTBf
Nh0IseY57cm5XaSzlUKahaqJo7hTYZY0XdtHRO4+33z1xuMk+izRTxDrFqa2BzvVSh0W5ST6Z725
z+N2aGXtj0NpxbqJZfVAs5eCckKnB3dJ3D34sUdMlIe80yDCNgtalh47z0bIm77PkkdT8SDs/ZGD
7vdQTCnXX5wTjOwy1TcnMrnTmE+ezQ2noh6Za23JoW5ejLZ/rw17AkCSlb7/ny6epY9CDUe6ASJD
mM6aM1FYJo0LlopUx2pL6boYBz6ea6y55GDnpS4PZ98NgWbqdWtWwpm1eBJ7GBYzqYKrK0/czBgx
IIDbpDKAmlVXxtM+aLwQZTWJm73uha/l5xk+jA3R6tgIguCUXg/LdZY7+ZTMUZTOTzBR64LVmU+G
sHRaMb42TvGPSm4NRFcQZW1NXVfm23a2tfsyfg+gYZUTAD9LBB826vIQpDF2Gc9OftiD7VhRHjjW
KLI5Mm8ul3JAJGN+OC974yhltwE87RLEas27BowiATcuic+4CbvpT9L9sfIBPUlm1M45+ngf6g6u
daEEx/jFLRysJuy5AXKq4bJyj58coSgGb9Pd9dIGxGrLMxPh1lwwsSb8AXWMyL9awGd363O625Y0
FoTwAwVbd+tFOfO+MYHmD6VbGol0cwa8aXQj8W/sVcNkfh9058iHBSobiD4FtkCeHI3Yzi0cMB0n
S6LwxaK28ZbwHYzQaPTvo21YIRlbZSbZ9CdIHh7G5zXKLqpwrFjqg8PPRs256L/J7pI2ZnzA6Pn0
71qyYqKJKPAtm0gDIKzIQybjs3nZRD2GVbLZxpI54S17E9ZNJ+LMBPaQPF+Yj28xSxe9T0+c+8j8
gkL5iwEa7J5fwA55Z1wKgZtG+ryfo7m4n2A/J4I3+Hx5EpowsrsVTAcvkbAOL35VxlmLjo0FCP+F
QaqNcnnIacVaNzwErkoY+NRxOdcUdhQsUV7tMFPSjWVtESXs08x/w6whYBMH/TC8iUuOv0lY9rdy
cm7rQIGoXBh5BjCAhs87zAVsLnfKFuoR3wRbi14b8SPO8vT4msF/e+a6Uth430j9HZqnr9qj7LfA
uTgkrgIyAvDr6Af6LU492MF8veAsSb4kQmQAlVmdfpTNcxqDywxHZLcFPHjcL//xNnx3lmZslg+x
ahPvHoua9c6jfDj4XwQkJQbsIlVIczVcNVgXg6hyPoMEBmQQU4/AMwOIjw2eyjmH7rwyoAK/ZPgl
j6csqfydfOnsW+CrBYECnHo6sETsCRb587UXRnytsVTO5cq/W776DM83LaYzPvKCazAqAPn/iYFL
AU68Zy+c34Kg7NB7LlpfgRwJ8fCpr2y36mDyScaJebAuh0BiWRj4W614fXFUgyuCdT2ht9RvCN99
I8NbB52mPURB7KpWz88gBocshRB2eSCbu38mgwidXZDLe9SZ29fW5O5toFW+NmESQ7j39EZtgHKW
2wxhBd5GnUfboiEGsL8wOUbjpvl7cim+CcdY1VT99KtvIKGgXLLCjepIqq0p33VkCt6SGNSg4bhl
gwJcZQklJJUSrjZJtZrE0hadt9MXRY+sLIzR+L+s5GD4roIeqEXjXrPytGaVCLqMWJsHePjgv1dO
xYCW11qmyUEPeGT9WJL3CMsdnhnd6eFppRmKyalHYwa3tKoLcWC+VkSCy1ux6sdOX2hmC9DtHwie
Y9JKUViLjkRMQAhyZs3QtgtNSGQbvW33Fv6ngd700PLXz2Tel5084SklKyJ0Qa5k13P+/XtJdnyg
F8fW9z4P6z2FlSmOT+PacrjQ77lS0TE3mHwCluib087ptz3crzxYKl3MQQQUrGAeVxL514TzQaJz
nygBR+O4h4G4EY4duI+WMgZR6MeVANrghqC6vEUlG2jUKKnn13G3b8RBGE0wQFrbAGQltbGRa4Ux
0ly8yCK/CEc4YgEJW6vsZ7AG7FiOvFZOWaaglNtSSQcTDSv7RIkdttDS8IsSYtrBkHf01JEC5mtb
JjQEj1RoATf7b1aR+QGqBuOKIdN2dWT0IOWsrMcxMKNWYkrNNsbKozwWGF89QDEiWTBd6i56SxhP
zwxsQHho81OD8uGuRq/yviOTnKKh7eUZeozTD/L3Y+zOT+rfbdQzDx2KREVMN9Dfkffh8xZNhWiO
XN4/y6ZieGdAw+RcPwstrU+Qwzy+EUFF0yxPQG5bNBics+zNXL8wslv6Xe8Egu1XJ/KKAoozfF+q
Qa9Y8XLgHImyEw4KBZuzjlJRij0RFohW4h8MGOjIlg1BelZ2IYQuH+oNg8K6vf7vONXPVbwFyyzw
EIl13HOH1We3R1foBhknD02PyOS8CBFh7gI47z534Y0tHKs5Rw7Oq87pB7LR4lUEivw+IdBpS/gT
z88CiF6xwbLP6g6f4MsrFTFkrtqglb2cNKHDVffsoUXAHi/B0BlpxQHeUJRED5vr6VJL/x79de2w
pYjJGrkac3yxsvo1tzmTAwwEI2AwNvP4xCYs4IHGG/0V+FSZHF0FO4FdlQkY5xQNsXik9fVUPino
5efNw9erO8SqjtXoqBpE6mmD0nd28pDjnhVeloZQpU84uB7LIeeLee27yL8aN6aLROMdiV5dgw27
egHis5un/rp8kOTDPMC4mutPekH4lvEWMH6tFIzYiBd0Z+etkP2F9XfA3VwVCE2hrJKxxVLBthlq
jTAaVH8gEQLJ65EXW40/Gh5wWnRK09+RAPldFwAaKd4zC+i0BEmYiZ9QPO6Dtoqwpu+Gr2uS3ddJ
Q+/tLliCA4H6yRHRODGOduE0TW0gI9Eu5GDBuprhH23QuA9PSvHdbtISwbeNs/omIe69V2uJeV2a
JkcNsUALDg5IZYUixlYrgNWcVXCddg2pLrh9ofRuB57pQ/dXW818bGhIiVa9sGfEg/x6S8Cphk/c
ecj7vHr7LjsNWl1IqGPbibVTMfymOapvrqNm0gccRrZFw+KDpe5V6Ew8rsqRk38+Wt1ur9sw/lhS
8wgHa9nUSizDFck51f6jjprzHPGlR6AQcoCNhLGvhX41CXs6VxVRT/APsCVWu/MquRVu/6h0cjcA
p5bhZ0sKszOwoUfmqaS9bEE+HDeMm+QxSwEalrhc7LKDkZ8QAOSYYcNH1IVqv28bdLlgIbm70oqW
Akcs8WBIOlKIwDj7HaKYdoZ6On5lYFwXghxGiIJD8swx1nqTghGxb0XpgWuIRFEQcJLdEf4VHzj9
Gvr+gWXO0IRQNLBtx8KM7XfqX0Z92UnobLzU8iew8q7nWA2IM9piW0qCX2FFYZ29oaMVKxHCP7PE
MLcE4KWd4mMg5lce2Zh7jouZ++iEqRCjmi7n9UUxlMMCxSNDzMxaOBwC0ZfoCuy02n9ymhRbtSHL
Ktz0VE7YzhK2HiJIqTfzWelcBafiSAahyJQyDAmOviriEKwNaoJR6s5I7LU/nIQLgzP6AF/9wdhS
XtQe/Di66eelxN0/ckzA4xH1WX+2lnfUYUPvG2I1bni4x/hE5dU6feftMKNojHY18BQw4o8MZ5j9
ylKSp9n717OZYHTb/YIJfjfIufr0IADscEWyskz1759oPmuX4IdNrwUFwyFfsFpM8hBQDV1sa/3z
k7cSCE54NLv9NaKZ9rjL4kuKZyw69hGpGn8m9xllY7oj1D9Kpa6ZK70Iy4eS43sXwNYylFhDuRli
1w44R2w9bLd6rH/jEdjhj9lwTUN4H8GluFWR0eKi9to95Ve5N+qM6aY0GzqxXU2qneFrvje1zXOa
fTE6s6as/1GRBRZTmlpQs+XlaAhBsxQCds9JtUAt5Zrtw/jRy2G+LfO1me7Y95EWG27TSHgUgR+k
6d+98fJQCMkDUKOuNpRk+U2PygA44lAIwTF4BJUZUgZmgz9e8djlZ0P+67vxnSHyyNGFxwU0GbJF
UEx7Fgb0YDbrERYtbdLGmooyDgaimjYwVKTaLuyzABp6MYvQBSY4EheEdHocYZGw4H9bbrhEkf/l
vcZ1GfrhGlgYOgWkMG9iIvJTnPr1OZpzAmiCO9MbiuUfsRGbu7uLycoDyMO9hwyC+vbvk1Mxc2+d
MVbB+eA6SLhAVvrciRXZLmesRcqESI4Xp5DXzhuw0EOt/IR7d5qZRQVzdhq+bjZpvFRk3Px59G3h
M5NKzwEvx1gTM3l3GSEiepNfmCK7AfPjpemlcExw8shCKE5FbW7DRRM6YLnA6JJOnVGc9+exiP4U
HdwpmtDeUk+K2+LpzRKIAe8ASwVl1Pbj2QZYLFCXvrzs9ivqNmxXNVSAo9N5odFSxjqrSoqyLbXw
15mT81yi+PMJQt2G5San163hV1Y8yhnoqkm+aPZpUJ6FGLjPW4VZaDZCsLIiVyX+MCcz4dgqQXcc
KlfXrueB2UzUOckpBjsmDwn9OL1TyMFlCyZ4ozgiuLOwcUjAbswITqZCEa3JAebJtzn7VFMtDgo2
jztjbgsgOBFKW1gbGgiDPActwQE4lZbAfJf+sGX9Giefh3ooLpzwpg862k2NOz09kVDjIw7uTIrg
OLQxQozsc934v7VaZH4qIvBvci6I4geZhF8PFKgsHaIrg7+TQ38ps5CQ2/Q3B52kUvxzmFvkwLSN
spCcDqOQS1rS8r9Fjp8AXMtCIQMm9q+On4cBPthWAaCamkmK2ZqklnxbpjL1YzYX2w6j3fdxFu5G
O164634ovjhU+mCh33KAw0lxrZBHfdUnKgKJZxi4oYqeNvW1RAXuFnsLXdEhf9oOSdDtupzPWuD+
kE/9VVLZ9Zvl9t+0W078fZmu/m0FkbzhTTHLBN3lfVQhKU0KaYfOaOnjBCOdafPRvUaS/XpAnXir
JWj7hd8mWXM+bOLoafteI097VzjAYSTVk5XYp+Py4Ur87XTyOaGhGpZBmRRZtpCqVKtENWlILB/K
jPt5B9lIKr97w7RoEaqTepaDrpiwHcgidMuFevd0OCfC0eMYG2DBtfJ0n1atS1m15gi6TKMFLGss
/4A/V3biIAtXY+V8V5aXN2xqLVxBm3IWNBfazxtsm6Cf/4+2gYB3/d/VY+yzDNCo8AaxTJwh1XKm
L/rOQ9hYHbXtiOXkBR6D3QTrmmdoTeKAb0qLiXzc/cE+Zp/43WL8MlEJhbHemnkkhAHwG/bOCd6R
R/Bj7N/nx5EJvMpfytUWt1X5ytLwE/hm92k/hHnla0OnqUfXWfaplThX53vmkdslyrJ23sSCB2G1
QaiBgrvY4VqrBi/Eizel3JmsD6rcvT37YxdPxE+v508tdTdXz+lR29ygCMaELW7vrKfH54WW1PIc
pPpXh/n0h9S8z4wMHOo2GZ6wqOCaRVG77cwwmNUAOHquxfoIJSxX7pnDYMD4VbyE2abs2m7L2l4c
wzUoX+Ge6sU4Hir50FzHqEjqMTABfpzd9MeWP8EAu3zVMZhWjQgAPKnzV/hhnNuSdJWS3So7FeLn
W8QzLEr08YAw7hlhCj9jDSs/ljnE/7HKl9U3QW3lwU6IzQDBRaMGrmaB+wY7krec1VajdcTmxD/4
hppP6xTLiDoaHzpVw3LtcOGLA2Z0AWphqDW9oP9DAg+8Ly9t4Zsx9MPz/j0pr6sJTtX3C3vnu3em
nMzaN6g1OOBhrrmdMnJ2Xh7UVrrO1/nKv+u5zQ0zLFwZFXwy6M01G8uLsPKS1+0BoPupyUzSusl/
fKPFUE0p2iH1SLNMpBqhlyBjBP4LjQydDd7Uies0zNWljmzqRcguNi6WANVw+5SXi6WQ8gRbCaUB
aMMnPWP4vQwSybJErs/4tGM1aRUXD3fQ+NBnNYSG55EGXm9RKF55Sp/ZtSUJpfLra482fPX6+kYC
L20Jbcg4NO15cVMcHRZVEAqlclIIgldI/tp90w1V3hdCQ0kOcFyr/URscvm28M2sxvI6qgiZfCl7
B6PWRO2I60eKJKqYdZiUDpr9WltJif2pMSC32JEoAmwe2Ui/JvJ4THaA2mlAUBjTorFJrGWij8LB
oxkoM7+eGMNZbAHQFStE+t0mycFYjZAxm7NeScNkmAfVJLbvIR6vje6rsOP35lg8/Kf6TENA/EFT
HpTzufdD5bt//WBNpzwUKN7FTRLkQJRGT93hYgEHmIlLnfza/5ZSrw6D2u48EdZO9LjMjUNzWhV7
nWsrM+dLFfQobizI+ZDwr7SmynrQw376jijXFtTg/1w2hCuZCP1UnmJzuyb41Y596ahNsiC1UbW4
LCevmWdK8Y+v93OGkJdWXPtO68XSjawCgiaa2mSKRCKNLhuRVeD6MFFiOZob+v1lL/sGVbXQR4AY
3a2eqQA034C+8uJ8WlOEXBDdxV/p6QY3TIIDyrUTp+z1fCISqQgdI/Y95HPrsRyfk/xwumI8zaKj
6JmhnEiztlTgI4tuTC5QHczxOK+ROFq6s6WtBZpDvrFyotJyQPbAUE4zvtrgtcgqsrtwmoXjJ/tZ
oaQQKChQVmNS1+dsMHM+EnygWQfq4MqOF3FkYwpL5GsOhA3J5Sfjhv+othWE83gRFQm4fCrjOBmv
k4zE91ZqKgTG33Sw9dF7SDnF6yyg+MXJSj4XbLyPdWPVKJ/rRPYQHtrRbuhkdIUrvsCTRITP2TAW
axRinctqSGy1HtZ+AbUphvbdBJOhxLHCfwYiatXHk0AXRFninbTv+zCMEaFGQG2d0DwAvqbHO57F
ZyR34zxwQWDh7Jv0Y5t/CnO+Zc+0/Fk2fJt30sF6OpR5ZtuCgT/MSPaXPfUO9Xi6rsgmGH2d8Dtf
RUOletMTYH7QZ7pGVCGxEPo7OFoTRuD+Az8tcjXZg9spn9CDWa6WuPWOmHTU3GCl+kZuBN4sLe5w
t3pf2z9zM9hGj5K6/gno3o2aSO6U5VsCz7iWOi3j8yySA5LaNE9C7YHl2oJA0VdYa1+uBNPq/w7R
8VglzOVKwG/FngXyZ1xXYIaG4fgVnM7wdw4DI8eUcKJjwOFi6GWY2/e8cj85JtrQ5opJtiEabyMA
PjZpGS8D57X9f0c8u73ddcQW2dPYdnwRAnMPONKeKEzcO6WPRy+oHuI71EgWQTfZDL3ane0hyh9X
srXBsAcDEgNB+CKLivNx5nBfBrak3LLOKdJttPifcn33gzaeEUT38vu2xs5gxTPhCMo8dVXzswTG
xKJeOJLp1ccBB/9C2fVZ4nqsC0tSTPJILkst5GkmwgmsNFIQ53vwn9MeVZfv/L2FIA6pjMbFa5tv
7b7rLUEkfRk8191MgHiHLft7rnnYxw+e+EfAM4hOdMq6vgILjUT8sQ7JDrP5Dr4+e2+M0L7WBGVp
4XXsT3AFl5Sszs/E8dN54H3zvLELtkzs0TtaIh0JFovUoxLo1gBtm9aS1PPD2TrpVAnM2cPtZvLV
CAHaU0UNK/vUEOH0EdThOKus2FaQjKWGvw/ygMLsUXXYlhbnzSw/KlYUlB+DEiy79hlueqhkVN2v
3LQ5fiAHJSzyo68n/HEcWTlHvJ9PWeqmEo2ke+MphyOhnK+sY3TcDphvtQmqMrBb2F0I2uhGTPaB
mv6pGf5kjcBF7sBLXGktwwOpGwwHzTGbcNSab6IMhHjdoamEYcinSmEWpgk3LR5RXquyfbvhJqTx
WnSUmJReBIB0SBM/lr6OvvqEpXeIAakbhRoTjTX5hewpgNSoatFZEe04+FpoKADSa5YtkJ8UvMu0
BQiBIhPtDFL6oIaRCaPRyPc6GQp5ZydJEz48N5TyTrhPP35RyS1/Qp1u8xr2eoxkphtjHSZ23Mkd
vrR/Yaw5q20dci1lZrkVQ84VeY+kQyjXWhTSAkr5jMHjcuxRL+999hDDk5EfdOh0nkdy5UWrWzk/
zcRcj9xS9ZdV7jejgF+RGopsGrJNolHhlwDIEarda50i8B/w0EUe7YgyMIh+QepUHXzNkysCenfC
qGnkAFmEJmt4xLc+2ufreWGkB86GqhOG6DcIEfyf4Wo2HqW1bNGsa1zgKs8sUfXu834NcAlDxeDI
1+0EbrIXlXB9EB427zXRzzsKO/IC7C+tQp+rNPfyqhHt0dhsz73N490sxemxJ0OsrYpKiH4dg5wD
ZTJI93+yd/u2lRBofnUwNEv2wOQl3FxThxivQAikWDRDWf7ZmQfp68G0hL/u9bisUn5Qi49LjOrm
kM7ppKpx/m5PIWv69iOqCVKMCnoJylP7abrQWs01mRLHQz24b3k0GDzPrszAKOxfsyucj9NAuwvH
+9nFNjzTxQ/AYSRo4g9iwEQjr9Kxh2qlU4gDSxucv+kDQoDwEPKWkMbAE4FoulD1G6QNzfM0NrOF
IVA0zxsHjAe/qZ/NxYsDUeMzEHJvr4PATZZ/Tc7ITpLUAJnYkxfHfOQDyK6aE+0sL8jw2TJg/DAB
gnZknNBzeYfywjtFriV3dLR9Dwg85PHASVREmXIdCEPqxLAAr56GmZRvysB6ae2AqvUnAfiTH9dz
cIVByfQhWafyBpVAfUpo987PNMkLylZhrW2O3DIvEJhiHnzZq6Hyke5wjqSLRFVQ4ZVoDGnT+7d3
g7H1os6C83nyK99CSASAD9+sAYf1GIBektKdKu1ql6RmfDQB+zm8nKfvO6uKPQf/2KNgo8kkh+dq
O4D9+RA7CXK5X+nwDa4dvAnrzGbzbTB2ZwR8Gd8ekVGQnin5HqwI059TUOppDhZ0FgJfcdMN3XNX
fCWYno2h7ZJb1Af8ykDvUMgpoTMvLWKMaCxNpbc1dohT0zlZsE2EJktbJFPMWzlgM2AiiN9fpMeX
BN8cG2lPv2c/FU8GpIl1fE+Wr39kJbkch49Y+amvFQP+Cem31PwoPSqtRUJPXk7/IcdWYLGbANvV
ZTaAW+h/IcpqqDuvyw33IksbH1/KVYFSKjfu3NTZmaHc6h+CnG1Ko+Qwkb8/qUYBfKtxC35rE4fw
e3A7HZpl+RDxfpi7Jl5EAyl5MjnTnyFeiX64H9zUW9n8NfnfFe4ODEs0RdEKcDVmFuAWEbhkoC1o
14NIvQzAymw2k9GW943K9sn7H74c73oHqGTYYKzzMp+pQ865zJzhhMrQNVATNjJln3Mi90kIOG1q
452JmMxV5klZkygIu/zRgca+kytXEXs6jG54KDpdxPZ2izkOW2NEd67ekuzoY7wf6SwWS+MMtJGG
9S3Yy+uKPYprtvF2cH4v0NryIv0onmNtLZxWTd/YHy34NMESwMejAtZcUDJrNdTZchuPh+blXAow
K/T/Vt/3Md76viF2yqSrHQInqby+NTqq0rlRIRG9ajSLdsvkD+ozOd9XVNBmCMyZZcXjFxoMPwkB
B0tB/ecuEOZPXAcFn+sUZnJTe9+zO34C50vsAFUlMpjjQfScsPdD+5tL4YCUxom6Kdpf80LRpaK8
/BKWrWkDtFeHJJwOw0XtqDHw53kCfaAwRguJPaHfnwUAOhwVcuv5rX3XfHAqUpUsKHGo0HN2Xdl6
AVjGSswxrsIjQxyExw9DCuJUZ+xgV7qWooD0CJ3BoC2ZkFYX3FkZtgwop037upEFu6N8hLsSJOaa
rHVRr8R4HeEHE8FOEBAaRAk7xtTJ8iXkeTU6L04ro8hu+nFbqtIk3dw11CbSdrpeVLad9Y13eug3
p4dlw0zcFglBssoiClykQJhr6N//Vn9XDFrpWV433ccX7GEXJEd8PCNP9jdtk/m24y4PTaE1AM8D
xNit2FLMC+Y3c+jo+PQfNUT0O1j7NObzVSXe4gr+EWy5RzZKJJLEsU/D7tzIDBji1H614y6+I3JV
RHTpfLQUEWCMWRYJzYC1TBIAYp5twxE98kna2NaZbCOkY9f+AgqeBXRFtAPFzlRYtkMylXavcARz
DUoFl6tT7tfXV5n+qVfbT8EfnqVGXRu08MRD3olOXtuE8cUoxdsN6NDhDt/iRWrn0R3Xeux1IvRY
UTGn0IxIbaYo0NNcGFALYJ1DO0YxXVlQg/DQYGCU4T0RBavrnW9eai8swmCuGOaR2W3DHZnYYrQB
voHh32SCvB+Ibh9D/JnVAQ18nV/qCizKGKFmGL5RRCgtVgRwCBvoCaO/3VWhpCAnix3bE52Qs5WL
QD8DJk+EZznd5Uvud0ARpZkoP9NjSnBA8lKjvgy96ZdysY2wa3Gqv4S65FlltPCSDqqY2fRvre8D
0TDJkQzOE+r/Fy2AlYqLi2NNohUVMbDL22xSNvNYzY84XYicM4fRAmBflMN3NX3EI3LF6Zf+RXuL
vg0jCJCV3vmIPVDG28/MdzfleQjNG6PuFcMl6obtS22rXDIiBEiN7Uaglg3dcfU3ivVGP55aUTSZ
fGUseBh7eS1dGN1CayPdbekCqPNn32d9ykmR29J2KU9+z2EHgVB57yIJGckB8fJmrH57eKL54z2R
OHW8YiYjF3HibaWfWTPyXtCk/a3hnJ/xEp46NHoHPZc4VzRZwDjOolx8tJsmQTkxjvFHT7naaTHk
yW9vmbE0UIsxEfzk/VtgeUW4mSaAMLqRRqgCLAj6jIccJWkOpwvEuiLbY3suSAaquRJRWOwF4BCX
AoCfWUDVEisoXq+rAwDsZMQxEOzdZcmo1V7vFRjxGyi2KxmOU39D3yDY3jNPHQV+H54k8twYE1Qr
qEqFv1flTUWFovpnLc0f5md6mojQ66UI6kDzVslqCvSuLktEl58GI7P5+m/3AAdCBWRZ0/lHV02K
49D4GBYzAdOHAlb2LZKv/zTs7HA8AiAxZq0URnJ0ANFSK0BZWf5bpx0h646KsOjPNxd4iKlGMZne
IRteRyiejyUg/EmOUeicsLkPrOUE7yk3KoBZgCNeMw7OWYD0eXTlyISf8IeNLQ+0Xz0IhW/JCG5t
k3gn6DZyeNTO+FQGaXavn+PtR1vyNjN8nN5PDcUxNN6yA3CrRsNlMupX3KbvrWjHLCCNpj/VD/yT
l1ToUCIkR0RPVkG/EoCaUdC3G5VwR4NX8WTgNOa+9NB9Pq8C4X6wMo/gQUenAyLLEIg+mvImzdmO
LU2MsGx4iaF/Vfg8+c7ZLp/jqky80S9jWy7qwBaVxc+1l+Px4AVXki3xlCYm9H7eh7Rwmu03Vbmp
tHftvy5RXoAI2ef5eJ1PNk9ljS2KuuNLqxkuq9nZSbO0rQ5aVljeSkVQYdiM2W4WtxXog1TJaQS4
GYc2eCvnQ+MI1Z9Dk9BDvY19maRoQb0nTm0FIFDTBCN3J0yJS6n8EVeRfAC7ttBmV9siDOM3QbTQ
AhBV80zG8By2LMK4vGWnTGvsx3k+Ki+ECohWOKJIctwoj3+8uCWZjgw9sKLLNnmTe8Lt3EnGkdPg
2BD7k5/w8a98zA0BcuQOYjLfSteXYst3V/H3et9y6fkDfXpNLTCmRM5eoDzosFgLdn9GOH8aIr0s
2Gob0e4NycHpn+U1jy4P2NhR9z49QaELdx/FlIeXC4bJoXdzHOjaloKUd5fX5Lv4ziVPRfVqnqD6
CM4S0uvhg/09xwWYmQYi7yAG9jnDiuVq5lVsfoOgYc88FEu8v/4AXQ8iyJm2kZ5dD5lBEZPBGmQE
uPDI9gLVJyxyEdT/k2ZJ3f420MJKQdTZPCFWbXsf0RjBN3wc+0KHZXyIN4/y+el4BFyuTC0AuCXZ
w8K0kGZv0nBxQ8moO8ad1UIcj7AnAkaK3ZkRuQGV2DoMt+d6yGzgWBUMIJXKGcekJI0Af7/gGvA+
VD4lPfRkWI2U1mF7hQH1YcSo3F25kZqcWi5lrThsX3zQuD16ppGiIuOAX1hh0AvmSIU7Y1fBsVuV
Lk3Y2kvlXocbblYbtGeCfB9CEhZXPcbdmeJSJTnT2K/IT1j9CjFmJ25AGJR6ExYU10SbTQBYN8DF
amWAmSQ722Bb33tFNYlOw/sGcYKC+NwlFOUquHx4ZXOk8XN0QZHtKcIQu6aUyAvWK2wncaqClFBY
/BkZZo43nytnWqP+VchT9JVw2W7NRR3d4vTqlavjv6GRKh/91QZ+MNz1U0TTJ3TojZO3rJVFhBVB
u3EuTrKMzj/wjtrG0srcdLQjgPJxQeNRL/yrpKxchzKcxhbu+IjX93Bzwd+TF8SSFzwTuBXmuxto
nrqbhSbbsUtuTkkzJECUaf7kZQ1Y3T4MbdOwaemAswIJHCl0tUeLaPlnVQNcF/iEvtZvtl8jnaH5
ROanw/+tUjuUaFhMEGtpYMRkbiPZlRByakoBTjOodPmdLOtAd/XFsmw2af8c2ye3gNGT8S7uTcDJ
PFK6H4PYUfVX5JDVZQbRRC5RpGefSN1yiNOfVucQGK4lixCGrTxwdwop/ryH7wbd2uhUi4ynZl/O
wscAopemkQMugnyTMG27lne0KYH1f28V/MA7STTpE+q4UEDlTkmUVROnxWZjSJt58pDmpB3W+5YE
Hc1f7WnM/w1rXe2VNKhLblGW5SsFNm6bFhnVtFty/aGZ1H3sGjanXAePNfoylTHJhxzE6d1CC2uG
9fQ4OaWuC8CckOesdqA8sts5B08iBs6ukjZuPhxSLycVj7nOl4ZD8ACjT/g2XS76F7CAEb0xvIyy
6LMVm/TrNXw8gixozy1KTr/og6g/80ugPyJ64xkJlb+xvYyHY9VKZZmpDnj3xvoz3Aw8dSna5NQZ
ZKd8t0L6t+0ksBsKXNjLhyCxPLQl/Z6GRi4+N0RBm72x2OKt140EwSpy2xOuKBRcVC+4jRh8kWTC
gi5uZLw1BVrDX+W74Pdkgn/7cGZabu4aNZEWlUYfNBfOH4XNsfuPulTJ0MCxhbfqN4fmKQLymycl
0pTRa4dbBCpFEuKXosJuiIeNO/YdFRQyz4p6useQEj3oUy+31MX4LKbED+neLJQsXfRLx9f0D7Yp
VH/aA0vT+CxL4gmPvBrqz86dAJAnP9ALQZAWrvReqe2wEkp5dNrHWqkB9k8j2qkHDl8bGue2tfp8
HfxkD+UEuy/x6I0Patee/TjifSKcYEhmq5zLRTBGThmiFaMBv5kg4dH1CtGexuh6AKqepfIzFuhR
hrjWfBXF2OyUtdY8v/0jKPOyLTRSWserwV8MPqkRmMpEzwUJrBhTK9s5f/3r3RZ0HiurnoUDI0NU
Wmgnjq5DJrp4jewNpgfUPjKpZnZUvjfXOObeeoY4WsY96hFfxnlXLgJz6+AUPvlnLUFsdr+Trklf
DgAcsOLPo+3duN7t13V78oko2/SwNliYi3qpfxrn+5A4/P1/42pPdZOjbQEYNZ4rUr3s1qce1SAv
+rycbO/XwPI8E/x3ZUStlwV6PkoOzb3Um6xrzMLP6AprlndFJjgN+Go2fJ7u7fIZrBcUAsszZ7Cr
AglQXK2HpiduxZTmr5jQfYFytBViH/JlS8XLlIUdQkMN+dQlvzJqMMpMsRb7V3ECzY8MHuDANvJA
BdlgOfrBrwc+RYAwhKyNkr2lm4S2HT9tqpjXsUQWriXDSUtzOUDvd/Bp5DUhCm3BujBFFMDRHP9o
kHHPxcmYLDU/PeBoTusMTnW6hyWbh5t1J/BiW+YvyPLk0Zwy3DHI/xQkcuBtd4buI6Yk9EE+khtH
9PPEdQR0dkIvEK2dEuKnSMK5ehYseqFv1wogGsbsLbtWuHJmlHPJ3FsHXmEFaxznl8jMyea0PQZ0
pt+GznKrWVuD9lQUMGnopJLDXKJ2FBL88HK7JuiOuQEtx/DZx/EZ2xrUS4Q6h+W3cXLqLCbKJ9hZ
whg7+Sj0wUwTvutL5JsHBaSeWpZYzauCKVbJgrCgPg/asFFm8DAvoCz9L27goGpXbLdhKs3XdOc1
ELwTlfmgL6hUAYW3wooBw8I6hfRpaxkqqyJg96oT1qr6n+bf9Sa8/g83mLUYHsoOJd5PtuIha9dK
N5lQZYgN5dl1RroJGqZ8ovZWnSmOJLd2dV6rWbEfEuKc8lj+bGz20/6UmGANPUtsAWOXarSW6vZK
VP7AeAUHuykUkCDpo7BAIaBR4vi2JaOPq3ISvkij8SuOaunueVipTaw1iXNSyJ8zJo6OYukVSiK6
Zlay9DWMwQroecWy5ShReytgW4YtRwqPF/fyC1auKuXwjlnThyWZGeGMgX5EWilknVABJo5XV88z
zAkGPES1oGpw6sHfayTPzx/y0doSESNZgXV9H7qjWp6NUM0xRYpVbCdQimpnWw/EET52yMF4Irr3
JnHMjS+KK1s+ywJOYkHutp8p3ZF1TTkkrAZ0Il2iKlWW+h+Jqq0zQ1YfxAtIBtc/CNDVO1ifErIu
A6mfJBsHs1sYtjJ35rpPoPJNqnoCWqedyLM6WFyRYsLaJWZqD1NoH9jtpVFD46qEMrnwcAjI9YKb
jEI2LmBTWtr8Yf0GP2BsQDFW7423TYXWsohNdn3DO9bwZVrL4X07x0ZX2VumSMl5Iz01BsrtnYeU
1Q14fc9visNOBwKMCj0UDgmCZyb9elpfcxR7kN+m3eIzyMbt/qg8s/PqDfWbZIReDq3ceZULHVrH
EBBHu6JIEDDvosX9+0nfalkKaIQYGiPTOncX7HUyRdqwOzv3UbHsEUvYQAx5f+THx5QwmlgK0AC+
/jVSv9/P/4rx3yHEof+qRI9iAEYGZeAVZpobFAJV+hbHIDSohFNvkxQEF2z1KCY+h53ALuPjYNzp
fEOLmiHXoKftlj7cKeFgT779iKMdH0GLukJSrk8eIgOuQoTgSI/h1wH8d6UEkFHR43zrHcaBAs68
LhgAyPN/KW+P4Or64tXPP1qQsP6+6mzVEbNi0AcfhLfTEdD9fGmI3wEIdMZMvhKJwQaEy0H1EtSJ
jRYAkVFgc9dw8w775xu8y3g3rbrAA8InlUW6rzuNV5TlClGnqgdUXL0GKJtIkJOn9Wu6teSoUOnW
IvgVC5hIPEzypDnkr9AqYb0KL4q2XZ1sZ+htVNT/0Cy5V/OY8bo4L2IRjqNB3N2DxJAcNvWCJqZ8
GT5i/9hv6XXXPc2dyrnU+PlF5z8xU9N/PAsC5o9ELJPQamO0iVHSPEV93v6+CzVfHdAcFVu3TZYJ
eDTMKHvCMtQASXrditU2gydblvnea3d5ijlkja/qawN5oxPi5R54DsNCq13NokjNCb+fM/ftYShE
NkUyYOhhM6QYZlrmAJfTSrj9BmJGUIwXQ6tELSMQbAWITl9yJm//YEMUxxUTmSJEppJBgKjafEN1
xUdiWzw085UOZBLYQ9+EtehhB7F37OdNbKeO/ZO2Mbz4622tkytIqqBXz+f9WRA8d6rUedT3vkNH
eiBke/T0R10gA0gNSv+5eq2ilYnnfCXdIyc2f1Xq3mBNMSnv9YXJ4cxNESX/llOtmDqK1V/wdZug
9TbNAHcPraJl0I6rNpNs9TBzGLeLWUf1WUmRiDy7mcA3PJCpweMZP/8j5Jn0AhdmGiebuoIMhTT9
VPkzSjgHrMS5zKoW/aQpLURs/R+ukHSZa/CnBKCzxrQw6h/km+tZd5jSDMNO1jSYdJOKjAjHWjTV
PeenaujOVRReuVjV1KC24MvAAyj34/TGfRT7S1tU5cTHHQ5ZOf43AAlCAH3HMpbbZQDIlUkgYPYY
mwCy9CuHvnfVwo9Ti6cUYF5KHACU1NmH/LcBp5/Kj8pE05HwJa0b9SY2mS0Y2H2V68VsGOLHXVz4
SNWvIU/wUUY3olONq3nO4E/PaZk9UeALg8G7bjHH/G1ntl2EqLsqcnLbJVg88V6r1H/yZZOh2mgT
5A9+DDLZdSna4G6M2IH0zrlTqRI7pWV3mVRe2ovQIiGXYAkiJiK6dqaizQCLKU7z9p6Ob6a+Eae1
IsZwnpUfX81K9YDC3Fnu26jSL8uUSiRF6Wl8jI9JLNNsNBS1elIJqcYykWDzWD8Syu1IHoiP3qVU
PAgfRFsVicg0MVNM2xF56AVuK6cJsn+CIhjGuhZz1F6xzVT567cXRpbmYDRzpyTrem/cUVqNQzY+
z135CrdhCTScHnVah2Zj+NwjkDrq7uBhxujWd+nF7sV64f885jiGEPFQChCq1AjooMaTUGXx04Xh
+voS6ATsr15LnQCumpYGccnYI2yAWNm1N6cKvXQUvjXbaEy+kmX1Nc/sx5QehXRfhtRtYdk6kNrx
WcZ8Tj3DM6ZvffsPuMlyzenGlI8HLk/93dAAyQPas3K7Rcc3VKTJKf36Wkpx+weJlIhX7Ga/0NkL
n7J6ZIQDj2ldMBOOC6puWNd5/kgbLlon68sHVavnHWH7GItRbJYd98EINPabsWie2VKRIvMESAma
4zKZip6aA1biy7n1VHZY4sEqaMKWA8i+j6nFukeTpe4twDem1pcQMW0sA8if/Se/fGd7hHSy2Pwh
fXLf5b8tkvmUcnYJ35hw3u6YaEFiWoOqrQiJgUy4LJHQbY0ZznWd4Alh62/eEY1wldZxN3IFOqkI
kbiueUJxe8gMUbI2pOci+HuouRxT2Iso4hlUb/A43d8FJeFUPvGvvUMdwiO3mRYIfEPgE9dU24+r
Y1Mng1zcHDXIc+2WYcLUMX59EgUceIw4cDREYBYK1aWn+nDldS6mVcieRC6BHFODn4dKwWxdlPWU
uXghUpwLOI47zuNy1w+yuEaDah68p98DWFtlyXhm+2uDQ5MoD19g/Y9CiNRX2U57qSIsqfyMsiT2
d79doRw03cqTXUHt1GDfSHgHFbK6i2mSIHjwtR98CJDacpNnamKDN5NrIWUkNTAvvGHkMh1XJS4N
1AkBNgW+2dPcnIpHaFF//zkwYxjpYc2w9xiYrcm8BeG8UOgdh/q6VJQhsDkO1oukf73WAjp71sAe
3G+uObyzORVB2pzfgP6Fwy2HiujoP24U3YkQt2CGeVFTcvsD6FM2p1KckdqOQHxJXgNK2SMVQIlt
udaPBqIK8JkCbg/7nFzlkWTtCOz8m5TS1vYxrUE475CKi2f1YCnjHLuV5s88hIrzel+Ey5XZ1cwo
pVf0SKaxpbA6De0iN5yX1YsELz7e2pAq50I8UN+uk5qANZm2iw/UJ6BeSEFnRJlGPnsiV0bLvU/4
6L5nnUfwjPsC8w5mIcVAy6n+dDhllV5o3yKKQ4kGkDs4jCrfLX+1D3voFjWw4gXjdrqDWDW9a4kY
GfXayhQUA5TTi6tWOEpLmR5+d+Y0uErqTG4CBQAQ5Yzt5IMZSzKb8dpzhWIdvRSOVWaTs+YLLnNJ
Xrq4Dy4YJqRaJntpw2G8ImCYclQzOJC/d2qhtzRyUU2BPwmjVPYz7iFFYR2dLfkox8OFFFDm4lMB
X9GrD+Esy+tsjqgp5CuWXeF2LpEL8PDqmhdSO1XmF5ZxpX3fP8wc9akJcLop7COrswBcoKjn24Np
/d189cTQjluZtDU6Yik1hMYEBKYK0SNmXaZ+xC8Wa5UmVRVCeDfSGV1BWDVwZX0c33KbsgdOlHJh
ISTQhHej+HlDBTXkFq1IyubPVmbEQLN+i3Sv3CVFlQeymWj0+0fbpNBMFA4R4j+E4fhojM4aKK6A
TgHN9tnNoB3Wwr0rF+asOfTSXj0JlpdCasIVeoGH/KRRwCA2+MXhT7jk6WtUdZDsRAs2OEoj/xey
TGbTcKgOi9epdNRGYfOsLSRW+RR6GIOPdSQkNPh+ZTbWLZrokbTXLbuuVp7EL+m9V3hMc69FNR1g
qkikW4RXH0mWBVM97FiO1dF41ltXn9VBdSVQnQAw2soNg5ZBVdgMFl5HXaBgBaQyzPca8+5Z/yPH
/vkGA2j0sDa/BTvV89mJ3X4E3ZslUV289eTe2Mqz4GXgzKHNJzPNuOtCWD/n6A/K1iFuPEoCDgHA
XEVociQ0yVwUktSk6Y8S/8WUfiBfKn0XyOUXdMVdmjLf2JBemJVB/onTfw+BMAQ1ZdbCTC2jWoxR
90+oqj6p4P0nBwccEZ5yH+4Dkm3geVQ44dIp645gCHYjByQof75eft4HR3RuSm8y3T8VgaWGBi2O
8BNM0K/cl+0YN/aUmcxFJZIXyhfcgZf+QIWShGILGZQHkGBUftI687VbpsZ/fN4FgaqMIoJJE7sa
KO0uhY1M6Lvtzb4vYJ2eArcid+LBeUz1eUh1JimEOfVU0Mf8mFJ8fdB/KCemGv1Z5Zd3U3hWQCUY
q+QAvgoNVeJpPwUduB8hz+zq2r3fCJhgRQ8IzO5wfhSAE1k0RQ43EATr6BBp4cxdy5McvSGUdjR7
FZakTU66eGrH+dV6thXAsP+VGg/BqGblu5FGzFrWlCochbXCN4W5r736SiEsSQ8osh9ETfENu2AU
zcZZRVQ3n4Em79aer5TA2pT/sum2Us/xTaSHyCFahUZ9LQzXwjCoil9m07YCgoFlQh0OSL47wGTE
s9N0Nmw9zgyC3XEruhN4wXK+xZPVI+Rpqkvssw8fBaOQ6lkhBhdiiiGJY8zlrPB/lPeIBKjtT3YE
hcgmOoaoFAwfu5tvd8+jOHo6I2PvVeBrENOw2Ht5/FKHEmvJiQheeFNqE9k+om4liLn24ak5Fynp
5vBPzNojoKBlSWhiB7BvvOCTkExjCmeEJsz6B2nKDijpa7R4kFnJpqU6wvs9TFbhh5xtkSBW1pnh
ZbQ6haSZse1Lt4r3Ui01syrgSaF5R0hyBn0AQt5XF7e5TjdDOpb3ZFV1Pi61yfXgKskbkFPikPK/
vDkALROyaAI/7lJvt1sMFc2jCc3rJsHc4Gu9PMl2K4J5LHYd0DLaiazYjuub8ghaZRZ8bT9xscqS
119xj+DppWgluAoJVCkmcdVhJs9U8u9VeLd6rOAQ2WxjBTTl/0tqx8mtpf36rgLmSMx5R5oGpPUV
XGEZlupLdRlVv3VexjrJFEnkUS9xFtZtq7qOS/O4jhV5hOcy0X/WD5OAc4+78NU9b51FGqLl/65k
ynvdqF7Uz7ej+mllGD7xEMDKQMj8MCzCXyFOPqCP3SGazTfOXpVamGEIN6dMsPBlAeYVxLWZiz1H
aR7LgznCOtbvfb9d19LgNJW1x852ShVBG6TZsdV8iSi/vKDLuVIjBTPyTcWI7qvft2WWbYH579Sc
bGZMQkHliCh0D+goaC6xnqwMmY/S/5E+fWM7OKanBXOq3kYU/iMYaA0d1IRh/eh7LmIaXeFvqN0R
Bu4/4P0EcJvJhG1lG0FtJz6mo8fjHnklvI0bLNnq/suB4P9Z+mVVr6r7DGTw/Q7t/FpeLrFHXo3n
J+dojazE6oWek2qQ+ulnDWZTgep5UGOJFWC+ivZJXfxFPkBEnt9oB8pTfOU9DPCeygY5C58cl2F1
d+GSNFpX/owOaSJrrOXqOVevS31EUqs2n3BpaPWK9yY/855JI99dw6FhXaV5csPUBbmRZ0zXTgsW
4QHWooUK/biD3y4lpJ1YcdsX7SmeLHilV8gUIKzIp2eWBPwTyhd+4n1+bhnvYefB6AROgZp0dq2B
zSRQb2agP3WBTP6UQDvjhGGOzn3rJjwx0Vx063KhLlj73NhWFL35L3xauXCcLC88czaARhBGNOo2
dgBAQyA2JOKtiBQmR8IaBe3qviFnYwfAfy0Ay3lzNN+vjzGQHS3IuHDvPu1vNLJuHWpL+QzAxcdv
neEcfiPD1uCiTbE6bi9I1Tfyed2C4cKXp8yVTAhphueSs+MPPZw7h0FHfIpvGbFMwXZ3Dy/2qUjc
2HY/JMeiApuHgtVJYOabIXpMRPcWKXbEeZ8P6WVFIE5QTOnakvNir5C5eaK9Qk0cz4pKeVhdmRdm
IbERS/cmzN5SXOYfJ5GrloUdttZK+pX5y1UzMRg/EUwjm/Zm1CxKdVtfx7IMnHQfZFtDJWkP7f/Z
W2LVNh5mPRf623dMuH6yHvQM5A13nK1GXKSbPOSu9aoKc63rasBLtDneC3qGMaZ7LLXfwr/aowfN
cmyfzj2KK6GYfjqricBmgGpt6ZTn0rzvRgnmNBMTZ1gdENPXaLKTj4piUgObrV8xtnlPdFlgCbhx
8UcTqiTtJnMen9xkSsbMpuR9BSdQ3zgymki5xYkC/SZkvdp6YCB43NEG4K1Ok1y1dUluQd+rCi8b
Ls4ISFMEJmeSSne0sxmlRcaaDq3sXy6WYsJmqRmsxYhIcmUf+koVik7FNiSbSzYKMjqZRhhlXfa5
JU8mPADQIfwdVuM1NHO3m4+6fv9sTiYrQTA9NyYUQoDSs/mEWJLoqEntI+MrOvUfrmOD7sTt0VFe
nzjhJop+iGq6Ifyef7m/AY2428bODpbisKDY0xCLXdnzs0qJhquK5K9pXmNDS6meQGl+5osfjr3g
ujQABc3Bsg/Temu2NOPcecsjH3aT2bIADtYraXHP/VfywPIN/IJWNSxJ0eIXEpm1upj2TnzpFIgv
P9oYQgJEK3OKjRamedXrvGRcgiQ/zFX+zlrSkqqpaSMfsra27II1JTrTE7DPvhmNy8ljNzv+/RSr
p+K5Fo9zk9lJgL/Py30wakcho/QT3EPerjjnTiYP6Yz2q4lUov9xzetrIiVtpYQCPiSGpWfYauDD
XIJAd2ga6Q5akiKUYJV+9WQjcooegbBHXjb1+on5wWpMGT23fNV1fiDfpjOu7iRTPVd0nhIU6L+2
fHAUcYy3u1OJH1JnPS6fDJiVBeqw7dNoE4Coq/nTYm7TSFnKG+JAk6tvPgAugmfgLZpEVHaJZgzX
Q6ECxFxwR2PMmlnMl1CaJU3z7v6nmEYuA5OxKuDOXmFdMa5vgrv8YtJEXLDlHnBuKHmiN8aZ0wPr
ogs3DGgZXI78A8yDXA0lWY9SrWjtn1/EAsu+B4Kz0AmmmLj/bGRenWI5V988f9Z9EvQ9HY0mh8XQ
Irza+7EH0CgKEgaKFVy5D9pLJA0I4HJ0B0HJRF7Yx09sg7ePDnGiWM305nPUKWlYrrg9G/DYNi0b
tYdTViw+X5h5u5yRFkQq9t0dNjy8oRHDm79Cc82M/bCTbEbeVDCl8cih0+5dQxVcDtvuKwL9E+D6
W0Lg59KOu8WZDLK5LBDK7SBcjqV7rP843bFt1xC0uCzmQCc7qS4Ar+D3F+kAEa9ikxPngqaSPqPw
5PW9iLIBsTzUr7RTwi+KJbiF3oX9HZjLzDtG1UrTtnp1p7h7m8OMTG7LPDzN2UPsT1UjFudraxwS
su53RvwqPc7ovDEJisCpvaRiz6m+ob4NVqU5g5UjkjWtX7DqBXYNpzkgnqUHKkyIozaaFu13wt3Q
m3xG8MEXXV2yTlZRWRA35yEG8A4mA/6v23TCvAGIBfgUSlRxnJVGXgnyjfLqMODcyYlAyfxYKa57
4k9YBit1bdP2S6naZbyyHIp6sk7vKk3lb6+YD9BjrBnlmI420Ux7tdm0zBPnY6Ty5miHWtH2r0le
tfk71RFYOJQ5kfW/Fk9DxEnl4YuxuWvmDdWdHm6lEyn00QIR9oipbMlbLbOVlVNrB0YCeUnOQbFV
v7OI+P+sLZZ0nCyh07WkDs7S1RuHRO1FJhwGcYY82XdNmeUPnebte6qN66a3EslLH+Wcmw4WlN/E
DNthm82psSfkXf94wnzzQwZniNJkjOkFZY1VUlNxSz9lEpMWVB52IGKu6s/ZAOnbR4bi0xX8pNv2
jDD01QU7qV7K91GxShPIfA5dmvumxlv7xnafpmhs3RGuxwQI4yoIw9FHmbTAcPKbvzdDqBP1K5Y2
aplGah+hUBkeykJ7vOlfx1cQ73haPqk8MglXVLQkRCLzSRL9dKMjbkjBWNlzcidrFjSF6jvAjJjb
jOrgbHnRlAuPWwibAMBsebn/nGcCtDTplFftbswNzCcn1hjlkKtrzOVqXburJwxnpK3ARbpeUf41
HfZZBzA9C2uxi+1KmivqBHdBEP71LAhurCRVvzPI+EVF1droSwOnisfeqX0htepxukbVQWucIwIm
jg1VDPMsBrKq9iVeIj/kJEX+svVDhYxPnXSTOA8Gi1gd+my2darKos0qgIBS2YVBR1cV2qbK+pBB
3bCPzIJFhW0itVSAdHEUMItphU9ugNoAlSgt17TUX/Ns+K2pLcF7wU6l33pfng3F4oGaf6Dwj/Mc
XClWLXCwT6w6OcUIWSySBSVsxTxBUD90Jvdmw1opk1YUKRPpUvHAa3l7ai1ssw6VyykCTyJKdNJu
Aok5pomlyRcxMMjCI3ShD5LcrRyrB2xaDJ9gQayQSxYYQxzK7RtKdRSgX4ht3tZx+gXKW+NJOQU6
x60HqvzV8Eu75E1cwtmLJWA+5DVFfKp1zcay0vgqXNdgKNIaGjELS6mTCAfhazkXSye+1F7wN56o
08FcEdpjIfBV31BYW71cMwZc0cLxKvZM+kooeLlrO+Deqouu8JbSAoi6Jpq528NEbUhWFJERCYoR
gZRTKkRjelcTteXRhh1ScudG56U1lwz3ePdcjWgyRF8qJv1iWK+JeBE1Bp+DG4AtLBMynf6fcXFB
m7JIVrBt2ZVashIWIZbo0s0Ts5a4GnJHp3OSEwcUlfQBB6QUMt/Alu2YhAmX/ecyS+cVHwjVBwS8
ADDvAJT9fpEKwAl1GhvPP1x2pik7Qv8ORvnzUcp7av8p9G5CLbpsmaVPhz6njU7+VC3UL0aKdEV0
H9O16ylVdDBvXcUGJkOuLSNnLR7Vkeo+mQVd9DJKCM0NK27Jq3dHMF+GDazErQMN6eC4Gd7Heayg
nUGHQJuJ6zygS/QbeXxVRUtacWsLnvAufErExxIseZ/rhDD+RPO5dBq6w4scrPMNlIyYuH6SApIu
5IQbsMYdqefld7xaWlFAryzyb0A6RQ1GZAlXF8G3uPl8Vw2ZbwLhIWz04q3a7hpLqFmlsMgKDOLv
cJhKVmZtD/xOg2A+GXLVkghK9PgNfH6A4MhxTM8ceJA8KndrYtQEnQmMlfKrOhrc7k7kUGCNguDr
50H8ytuKcP1HFd9YBS00lpcutld6r+duNXt6CAX5ejnumihbD7vng70SQX3v2b8GtqnR+8rIURyX
OS3ZZnhJ1n+p6qctfZXZsgMRw+s/Wq5tggDfSyk0hzhQq/VoEKRnUwmnIqchKEk1J3UFGCAqDxrW
1ET5uoT+0ZWT+FVzjfhLfuZSMOa0Pw4SLFhPLuhMOxAKSsCnhpZRRX+BIzwk8AU4Ab5RTU+xkX4w
pYkCE25tDEtK/aVaHQSvkrOcaLexqIyCy7HrV6DFUmDqUGTWNhCqbbcgMXNMLpOqv65aDNsjKWV1
fSpHacRnsm6p9ErjeNl4ftQsNR9D2FMPKlO4CkFGp8C91CDqw0XbkG5m29B57bSIbujlD4TxWl5R
P/ETGf5uKARXuCfuJnIQA7XrSTdire2HqgG8aTmrHrCBunPWeJozqALyTy13SzdZpZesVByr3cnf
19PcXmpU6+AMLaUIE+IZZJIJfYs5E0QJANTSy2CUKmaxXv6jtCjsyv72LhHbfGUBheJ67CMw3+C8
EBYB8OYY4LHhrDWqQegskcziLjf29W8hWsRtBioO4VrB4slTT5/f6waGOsDmqcNdM3s4v9s117hT
H88AF714Vma8bLCdbvhRD153e+4TFToBMI89zOp9IhD0D8q1KSvMbxHIWnjer3Aw9jtIy3PXKltI
SPpYADdd/Yxo4DksfyjeKkGdOQJYtdAx/nLMU0dE6PCgJwNBQufcZ2Asfaxt+te97eVIJiO8XUe8
jCYd23U+14nbQobf2CEK9ElTByGC+Qy2tMMP1ck4LYah0OpaMOo0S3XHNHvGjC2DdqvakkKLkhHJ
640ZnxvhiQoQYgDeS9H5fzKkZhNkEocxRUjkfuGW+4Bpik8V7xDfyUFla3hlzahILnf0CU/J5vjG
m/47E5NcIBRkvccOuHFa27L7FBf8GDvORDWRH6Xwi4Ddh7DFOxQWjKQCcZjq7QTl0fe0WJCHyPwA
ODw6eGrov2U/YKDrgqto5fBLVJ+JSmjZf0PuOJsTtTlIrFPhZ8ePjq1uXoiUEIAQ870crMuKHGOO
Fo2RwcH8rOAyS47DKuwqvTNy9bo7xCKmqxDCQLhgZ/EdCMSMXJf/hiHx3YeGwnm3/vmJOW2Grtdn
55wuIRDgDVj3RqDMi6crfIGrb4dEr+6EgJsqhZUTZWAAOakpWlmDVxI5jlqfhqAujebzfNW5Q4Pb
hJXOs7QhrdqlScPHg+HQGjRsuq9T60Mwnz7290x4tlDAvZfvkQHRuXdfjdYPUu+Myw92LTAzDP1z
tH0Vj+OUpURaUdHnTqO6EY2QlUhFo1MPRP0DX4xQCHu9MUPSkUcOTVUoESt2jsbXqURlquf8ctbG
lZ/q8iwxd9S0YQdckxsu/WK03n4MJuiU6OMtJlcBJ2Oo6oTyEDdXL5Z9qs37CpIm1XyXqrflCKNG
9q+JgEz2cWK6t2UCnqry72TWXJ0UvEjPDwE1NdnpmCa0knDKAXWGnWdgb0ixc3KroBD63Gt3c4vw
lEjfwa6mAySFOg+DOey3xoIZnhAmdvmvp4xW3naAT8IHpGiAD5Bshg7Dg9O0gjUIMkIhL5sR9A4c
CK0nUe50mi0NMmAMb4gwXaPUfm344BLMDUptkxpsCAkKNmUDphtPD+bp2+CklS2YD+2DosasDNtH
4AezXF6G2wVLWXVMc9r1mkh/N9+fqu0JDw4RWZx22fxuWcwYmxzXz3B1CC4PuDc4wuDtnWDN9A8B
gwLXzYucdJwa0ktnqeV6ieCTiLASyFzaKJp6V87t4KfLrPbaFxWCGhUD/2FBBOpYpRA1GF5I8hpL
ODhc3QW7utI0Aj17GYpM3mO71B76+SIP+uCKd44jnywRRuCPbZ57vEnQqzbK4U0g3mwpvgZisVWq
lMjwvdK/M5mUF7KnMBdx/UNLTbA82ZInxM6I5RdAh8jTsGyytvjRtnT7YeoxXX0+CZszU2LfH8vy
puz6pQBIiBAMTJA8QwJoyzwfCUeOZGf97pq7dpvxUkgduXNUvgBR2rqxdM8VC84IMlT94cqjlt25
/b4GtroZknS1BJMyhmDpVcnqIeXgSNJhtW0UWd+ICfQZqlj5hoouimzLZhbX2016mLUOaBdw/g5y
4hpHnzahpRPaEKUfmTC6m5t30gkLON+aVaJwkgMkigotrs0D+dio/lgbziqWXpfKFVa+TVzRpGfy
adq/ZI78MsigH2+boN4dTjX86UsCAy81roWC9YUKQOuiCqL43IfPd4H8RUKDtfYJUdAVEAClSqhC
SZmJda8kYqsdRb9Rl2GiqpFYWsQ+VN+lntOBl56qig6dcz60IOR0vVB2wEbp3T1dkqYy/kXl/CW5
gBij2gsDcYC+1boGBjoo2hdX2bn1fn9p5KwMcdJ2ztlg/GtF0rbbROqI6EZbpF3xkxUtr/KympNY
CgcE5NXp201y8+I6iqmLuzTCdULFKRr2YrM9dvNrQHc9rwFBVFTZCs41VehcXrsvh9a8WvjzSWTi
1kmVDwXfFCdElmPUVeBU7KYkeDoL0Z+U8h7DGPiCFGpJ7hZsPZPT++yBg0vrVkIISUED/DG4wPQf
yvRvh2JZ8zV9I04NAx0fgS+QxoZkv1J53jmWPJzjIEaAXtBTraDlscDrYyRIKNiZC5ii3AKDzjkv
tsSXY1tUfYsoLHDDuFnYL/lNRtCKH6WCSWUMkqFOfxlW6iVTmJhmv9+RoBG1KKTrjvgg/q3uGsw1
xxdoxDKVEwCtCbzWkTwTCEbyS18pqmUxrpA6gQg6AiuurccbZtPdUuafLJVPPGtC9j3R4t7wfh4c
vtu3iqppzTBSlS4sOSNtlUiyexDrogv9U0EEeV8vATWFwhjYq4oIILRPCqAcZO26JkkY96a438oZ
qi5mz+dXHl7tL5vKy4TaXQ6R+1iqcHIXT3e+XRFmqqqiltvL4JrDHW3++afAisijT0zMsQ4BYvuT
meh/timVDqM2RAVDHWxvBQ/gLmmjxVvPCDTItpHs+369gEBKvrvoYlAYksqYZlqyke68ct1K0YqQ
f6a3fwr6/vahgBw4uvTVWkFXngyFOrW+g1s0qPYF0PArrArjklGzdQf5GGtmRdauGI9hBAKM98Bz
4FJieERmMNlYNZ9HI9eVb1VrL4Te73xvSz7gcPe9iMfFfbeXQ7i1tceqGA5Fc9cvJZ2NhY01VEEp
qs5X3u1gHlPh0gFf5hTjFBy7V3kTk+f6ckO7Zug4vpK1arp4tMp1AjjcWQaA3tkRKcO1X8q5PNHQ
UpMBwCRo35IqODmJZlrylKSKlQv5erVlQYh9Tl3ulXwF7Y0AAl7vXCETZcnSgV/6gJb+INJs+Xyb
K/CKKUoYSxZozAN0zsDCyyqUehKf2ntFGU2xnE+GyiKpi64tSZM88DdiFnngj+McOceQ4SDBRxJr
03fREJ9cG4D6pYJNmi3Wxj9J4VneiXs22d/4VUN4nxzNTqeBZLaznKJPEOAqwBk/aNz2PdzgQ2Zn
UFkS1XGgok02O9b4mECj2ugMbtg2Ot076v4BvvDYi8gG+RCC6xNEzQQQbNvnLejlo4/B9R0YOSMK
+BA/DTd3MQWKm3NbPN71Aumgia/5qPU0mrEzm6x6GyWSpHyvls7JHRstJwtxxPHuvwkBGTSUPH0m
81PUQ4qpticA72O09ck9mvjdCu3aPvJke1FsGWE362D0CkMrrQwWP1awiOsVTksTJDNvb3cdVyBf
PXVAmvESBOoTg9YgzfJSW3VVnkEmRPX7CSKLcCWxyCjyPnE5V6eh4yARzgzbzAkBHySyWMKbm08H
hbybaodVeEuyBMiBxQIQUohQugRIBgmNATQzn+Jz0dVbbyyW5J0n+SegWFCRXYI2mUeLrUnOFLIm
i0clgFvYe61QRbcZWHt+9Lri2RmaEjKVzClze7SRotdWM3tlMhkoAHZqsMpjT+IQpGBm3DwRh9nK
VIHMbicSlal3jgnrtgeyfUP01pAh6SJDZINoQl8unkH3L9fwYuVatzjoDbhb0eIPSTurDcMPTSDK
ehoNWmQzQxZAVrxFtfYZHMVYnvUhOC8Lst2EhkNW/9riHm2K7wSFPMuqE8bG+YEZQCc67WMO+MPa
CLCw/DasLZUBRvUwmbSes3DWnKk3iPdt/ToGqjAiLHERQH7SnF4DFilO6G4/ZZDCZZvKOhkUUmQ2
tNEbkxpjIp4VUYE0pv8L0ENT34GN3QDgqgtaLGE+LoN37yrfK5gjq7aj66ysJQrLSKs2x74t+35E
7LzU1rMSll6mJyFSvwFJenAZJ0MCH15H7swyGD/jpxRvdTM0LiZS6n2OVFGQOJyd2yl8cNeo3Tjv
7r6mZLjS58HBnsdPcHk5NLYHZc11/SsqoW5RUkJYiLa1JLrnlADPWcIiM/o666tAzn8s2He7h/vv
G2hNsHCxi4dQrfWroBYKiZ5+z60JIoDD9p6EOJNAyE1/k/aPHwouhP9reoUaznwMvmhiHSL9cKVm
QltuFP0EGQBNpU0qppOXULn5IUDeVWVXUg8tHmO4lbee4nzLjpAHUbfLJt1d+AzJnP91+KQLT7YL
kmXcLdjvZAgsm5lT2JOr9Y9HgRSoVabKgVSl/IksTNsUGz9eIciD8egTRd5g5KJUZzLGvK9eGleU
wfhBiBax8vsiCo3yKlcQB/LbC7njUW1tn56AmAgbM7cgb27cv7iZdV1UDx5TXkdiXxPERkCHiDJA
+5ezIbiDlisLrJpeauuSzvkY4ULLVJPuuZ6VlfxqDSn0moRZni2+9jpqoY1epeZ/IE8AOo1NF8ml
WsKP2sfiduhB6nDWeFkTIab+/4SQyw/5M5AT6Z6ZbkyuB4uMEhCEz45akTLwhqstd4MD+tbyJhjj
7dOzPalZ0G3S2BqmvMp7P3iQEeHMibafjqgil5DvDaok6EvIiz1Ldx4OUUG17ivTE+A21hvZe3Ye
/rCownZzQEM/obEpFd8bT8qNmM4FktsY0cJWiD5gZ8MqGA2t/SDWNpufOIAda+eiepnp/aWqcY2A
RCRIYiPvW5kZK3Bm/8T/Zr1jYeEsBYj1C7uu58UTUbE6eseK1JtUtL6n6PhYp4c/si0RX+FNXeNl
gTtoHeWuV9ZvQu+7cUbDwIbrt7CvjNqton3SijpejFi6NwKoTtvNiis2KZub6GaQsAHhqIxQAqTh
LXYz2f8CKxapPokuyTaLMzWp9Zhw/HRePSE8nP5/g//oo893BPYjCKo4ZhwxUeUiKm8/n5Cj1d57
0Qo8l+z+YL7NTpVfSNR9fNhzO5SxekqUR4F3ivXHLjKi8txRz+FYCwG2cAqlAzPNfxLjdDmvMLQ0
opSQ5iyM6fOT0yvUl4DtrUefbqA9szEXTlsZIJxLhXocMzN/5iUlgrsGiBlhVee01PTLFepRLJIR
tU3Xcr5+Lx4MlOWjzmOzH4ze/IUmH875b3pyZ4rZ/zhkrNwgHFiP6e+6LHyMXElDIqpn8mLn+j7N
BrgerWyesX0Qoi8vBvTts6IxQ8s5wl4bJHu03ylLftOqAslgA/Vnj08HDuG0ZakQOdpq6zEFnFiZ
YMLJHiFwjr8A325Bo9BLBUI8d6aLunfExjMVunmnzxBNAuMFFc29Sns3aLaZjHOQJmT81ZrYQD9R
NEOir5pQJhMyql1T6iwqt0kuFDwb9IlpqsOL5WUT5E1tc/sFkqQHOPyL1BG0aw4Q3uOLz0l0jmfC
sQ5s4K4UXoK3yJNzCDaMOiTvIp20NBMn5di/vtXiUtUzkrsK0bmxQDzXm8CXv4VuV+nCl/sQdE+Q
4BnSM1qwdnnsSk8arg6F2Jh9nIIGlHTUXhi0FOepDPTbsFMv6ijpgefE99Mm2sIRrVaMywJeg8xF
vnrs3QTtXl4L4GJFX4QJGQo5SEZm80nOxgrfkdw6n0ybzbkT+DFkEkOMgEU2pMYGcU6S59ERcZmd
IsFUlQndcrtE1TICf6knEE1fgK4kUEzREMx8HdWSscBD6KKcVkll0HnyMaaHUFyU4oZG86HTcKUj
HyIencfkIa4kAGgrRat1kh2wMnR4/6rVFVq6rYbYuqlCqw6RUXEzje2liEbLI/HntHVY++1DFyLw
xt51Sm8Wfq5AtcYbpIR/k6BxETe3STBdVKGRT55w4aA4ZOcstk6x7+kf7MUSqLWGGjBq6MGmcmz8
t0Sey428wuALSnytJr7eohi5EfIzkUV8RfbYXa9l48Rokyo5qh3ZtRptbwvxx7XDXrpCgYwgCz2B
w6MVTQtVDPebo5W2NDi3dYHwMvnmySoLUtxkpnm0PteJCxlktC3qwpP2xEbIBDSrE3pTng/99Y+3
mAdsnEyQcFz8pNy3v1P5MCc1L/5LI2nDMidI3dw1WxgY3T4WtbYeBrC8Gwbxdj+N9BjPQDi+BkD/
Lamdp1x3nJ0SsCMpVfMljzNu7ayID9h4LRVkVNo9Ffrh6col2caPhaUXHH1OQjhgzbStrsZqUNkX
c7ydEeOq2P/NthI7bEzvF8WNOQYGDOc2RGuvYL7HunYwcg3a7iWY+Yru6IrVPiyK1riP5yG/ua3T
7mXrvIIpPJ6/jDpHx/Sy+UYkP4Z257ej4Yf1/7XOwJvmPzT+wSbrTvM9+e6P72R6Vb2GmjACGCjM
fu/bo3MEW9eFS67zvLF0XtX7kOCrm8cwgOMsO10CtfEhLpLFCQtC8uXMYiqs39sVGVQGIfhZOU4t
s8YFCzBw8i7hn2ryfKdZtaDITfflvkLWXRUC53JbOSFCMDa1jmp3CMR7is6HDngRHjKkbW9Pit2m
WuZ7XQ7SxbibU+AYanQuZ09z++f4FUULvBU0t6M25M4UqR1Ub5f1z0gH1HX+YeSyto9kcummrHS6
/XHi0RaT+cugXGLON0qWKSt9Ri+SAQNLuHj8dWi7hN3hx7MhJ4SPpORdi+ZVpK991x/Z9nbHdiDa
sljwqzotKI09vlaTSNcLy3vc4td8XE3Zid6etV1Joj25RDLi2RlyzWKiEk46j3umIHW+TDn0CUY2
qFTVx2j0IzJD6VqmuQ4K3fBKQFORyzqJwMPbT+yRFE50Sqs0cAvUVDkax4RyQJ71wG8WfI/2tG/1
IB0PfYEv2oU5jUTHAIjkyXNIzP/RkAhHQrBK50tiI8jwGnFp/MfS2rNp+ZBK7qKaKTOeeKjn3myx
bH7mYiuyOxgYhhu7pHHPt5FfXLfda7u70w6EsB+Yd64DpwPoRWjukso+uvtv4T9uF4cvGdc7EN2z
nFlCIM4bwVJonaqKDrGCvj3DpsrmJhuhlvgq9dL++c81vMJqYsiTDa6JSOECZqBjjqKGQcYDObtX
Ea5hLz0HBq/DV9VKqBdOe/b7w004D9eKzYh2+x23LITHoW5Ts9JHEIOoeDytOQapfPC8CFTogL5V
dT7Qv9qEltCcYCKrH0NNn7twEBrp9RdTWhgGEQSav+0vrg3Q+A7KTlh79s+T2bsqVgsk1LxmZ3/z
WT13u9fcILiQH2jW9ld6YJx7rcVj3cJauwlPgXb1qVuhLqFoH0gIuHS4GiGmYsZ8tuIRhdTDK18M
cTCJOjT19c2NUQ8cUkBJ3+k/GViv2B7hxmILrAEkdfwVJOpcRcCv7FW6If/Puf8K2SwBCv+uYur7
pXjVXaNIKF4PaHCsjeY1EYdUnnO+1yiyHHkQInObvaIt7f1j0Hg6wBJ/h59PuJTkNiqWp9dWH+z7
kmYbYnqsIZKlUxVJtuSz2AQQiZrbCEjzqxszoDQ6OzFla05rjQF9jvocuQHh1URhBs3hVfHe41Vc
Z8imH6GePkEcfbSO6wabSL24OMUVue/X0o+bVlcOekw70oesGFUwTYrNP28kvw0M/gjOHSb50TRC
SiVCYAQgjKJ/y465jrjQbeH2uqGTOqhYZbipAdHMv+NGcYafLEaY2uUMTwm4420dIOHBzKRC3GIQ
hsm6Ru9mt+oHr5qWZqCQGvuQgbe8ox1Z5HcTPLrsfajEZJQbx6ILkpp+cbUB/iYFiVSo5HUq2n8L
sH1rynOPUvg/CbNxwmRQJyKmTU/VX7fvXXh/kQ4mwTAe0U1CJhUA6e8/1xZB+27OWeIoqoqQ8d33
7X1x3eFCBrTEwmTrJK7+bY++4Vvg9K0JXhh/BCcHD4gWYDVBOgcwGDJ1LXJ25LpPHhDjQZ4Poh6f
+J5aFiWYNeIKRRNWBwicppfpEK2APBfsWOVC9MUYVSsyPRAAK8m8fK5yorvLIK/ASQOI8sGAUH+H
ZKKu74e+F/WIVee8TVpJM6jRClG9yh8KOZFrOhCRYgxr+JS9AJs86hEpID8aPOB+pdnO/8MTcE28
6jlCg9OJbYDRi77AdI+8QMJsdRNCnF5xrpYZ1S5TLGgx9pkFhd4sqrRHXTNKa+W4v4Dgz2UEoPaf
xzBgn+2uDNYjzTda1eN7vLQocXAS8UMjMpMyOT/dwX6kk6fjIPecJoeHxnCQtnV2f7k2kdyufOBw
i8dAZ5bBOHsUhkFQhtCaqffLHUQ6Rd262wnGVY4XOhfGK5p5xC88RB5HcdgSu9HTLyvhbYOxJbWo
59MMD/xqOCJksWT1SmDYwqgyeT6fu0IqxcHE6kaxZGCDiyxcIsrWpoXCQ8psc6Le51T7Wd2qRpo6
Ug6otwGaWyWNyT9Yq8bJ1Sy3qulmhCHeUdB2Puw6Gr1jkCk6iJHR34fZWDlTFqgUjg+RA4tCEI30
hWK0CN8I1JpL6bjkiuJUNwvoO1IWBFYjWZHNG1NfMH3AWZzo+FZmNlJmOvMhFUX9n5YdyUrtd7Br
4p06ndruBs1DE1uvnPq/N3YTmPIboTCZL3m76vhqU5QCrg8l6otzCB3stkX7SE6CwrLtjVA1AFtx
8PWHeGU9DQJoHaRLHPgWEgk2Cc/SU09qU3eWMSxoDeX6h9fgpTf+DjmznG1zQGpQ362+El1FuHjS
u9ZeBz5voUXHCiE61DNAMbzKY/QWQEgRx2C57JrGYDrvaD0/x81Sv2SfOD2blgQMcZiUSwjTekR3
t+fcwQK4sNW90X7JKxS2I8CX1S4oB4rTGYSFCI0nXpI6wRPKb678pt/vO9UO5l9La8TBHrH5ft8g
1hAh3kD08q3+Ub9GpwvT8wBoRax/J7EJfsGzJUcxqODRtsA+RxoK77gZTSOZD7GzR46kwKWgS1/s
lA//lEiAMNVXALKguYuGtfV7e+KASPpUDULp5kJeNlYZH/CvPb5a9Ekyfwkms3nE+52hwc5x210G
brdm/whJh0QTkuvB1gEib8BqJxYb9gUKCfyc3hrHHq262D+Fwk5Z9lKPTKjox/j1tSxmyQLpnySq
AQQpkic9ZGYbhqEArgvjAGrS4QUulHLhHHsDinlT10QtMQZXTTKJzWlPWMrDJKopYKFl3kd3DcIB
jGrxtbAG7cL4mfLf4rRCX9pntctI1ydY/nxhhLZmfaUyGQBAOH7N31EBl08rjwJQW4evTvQgTXB1
dtsBVdM2FKYIM7wRKFk6T1NyNyIEZ3ekUvssxyGYn+3W+6VSa+96N6hAWRX0HepTYuw3im2BMQqy
EnD762yyD4jTvLHvNfSg3cUlJ1WMEvDPyL48R0p1tpnPJXjjJ02upSZHhVcaXDIrqg6EsH1oBFDe
Sipc7k00ERjR6Evhq+QUlw3Wi+LbCerosJCBJn6Pjr6g0u3PBl1UdfWZ8+j1V3v8ayacuwRZFj5R
fY5uOKPYBeZp9VE7BHLobO1TadD8uDrcqPG3+gjT7mJUM18M1RI1B35xn5iCB/5QsqjG+cHP3IAS
Vnywe+qrmO77vWKykCTeuJx0QuksgwDDmEswYzG+EIb7Jyh9QUsxnwU1TE5K7lU/CIhYHuUFEUCZ
K66Sxj0axgUimBmty417zaQtA7Q/rjmkRM/867eLjCHBd1ed1igpS1XLmEMYkIMoYJQAVCOJGRGZ
IIf7tLmi4ZBWtjXKD1EaSZzZ37zOPzOhE7dhVUPr8+AQRXo4OTgIaVgzelpCB+0RVqsqLmQszduB
zw7JP2j0Kd1pZY1aFwT2VEEVXWOOPNdLDcgCqfJ6PvUSuDcENW+3gdS/9DzQ8th8EK/GnwcTGNYm
cf/4IIrs0wDoFS5gwU/FA4JwVOX6vSlAj4bBiIILWWKbLv6WKvjyvlzsYX6bpYZqOYoTf7A9hU2W
XMkxiUm6RT7iMzoL5vR7787etLdZhyfbBRe+n6BOm9wYd+QIVJcTJUc3N+AA87vK+chDKdlYolzW
xbtlSUhf2ss9Hd8BcHPkgdViUmauUgiiiKRpaaocNs4kBXYGPZMFaDB9BZUpnZjXkazctZW+wN+9
1ZXAEyhLBkaUtywP6NRQGpVxa2pLUgbquxg7z0TIniuMYbjE5hZqu3BJSa24qOtiHJV0FUxmemIj
SYpuG9MY4WjygcjBuKAVD9NVYjPfetopdaIXa9wBzsClEJVYRedy7iDsZDyo4liVSc6/SEbEEiAK
Jc8wq3/ktpYDIZWytnKU/aYPpnhQoox+Vr//CHNDdwK4LVxghgSgxcGQMA8bWuvVRbLt7J5dRX2M
j/6xaZKIVG0V5QeJNIsWtT1+rLeoPDyPhmEHCLrXPr7GGDBcbGIU34lST4vIJOAqgt9H8WSNd+UC
y6zzNLWAMfJhehF8fWjStON/O3AvaPYLrRVpvvvivQNjUK3jVYxKL6ht6AANTu0jmQ8IcQdAf8OK
FuwPUtbdEX0UZpfO1JVL2FETKbt8QtgRAeFhpG2zX72b9p+svr6MnwRAcEOfcpp+sqe+qdvUNN03
DojrUJ1K8iwyawIm9zJdTq1ZgyPDoDSmKOpJZKYQGZ1HmfKPHaH3fW/4GCdotTl1h1UbVKGD07Ms
5x68PDemVLL2M3fUOm5Q5Vk7PAuae5R5EV1FdYe5rUqcMh8FwGrvMP5RHnqvEbCgvRyAO7htdFAb
STsraTWV3M1VKBaLB9LlBPW/R0n+W8tVu+VVAaXqUeyNtCMpicDM6A3R5fISCAF0MtNbm9a8w9ZO
mC/ZGYfx4214Y31qnw6hLkWpzaZAvHCqvOhU9lDeKWJNIVdAIoJIsxuKEyuorD4wvqcDODM8m/OL
rhF0Sg2ZGJsiDjbpknjAyL0f63g6vgHlrzEenRUXgafOB+OPdEsRYRq05oaQZJ4knppEHSCZxipQ
Chj+eloLzQmBt6nW0gOjfCtpw7W0x4rADhQXBhmGsT2EYBlBsv/KqBmQwWlj5S1Xe99Cell0bUgS
ubWTYXi2glvvtjutk6DapmYB9srySIHb2bbuKM1cq1u4dAqmGwskULil7YJ1nyxrqUfH6+Lwmw/A
OlqK83qY8bGTPMpKxSyI1ts/QmcQFDF3mX86l1Rpp1mQ22gs6XwjuSktQt1vWn/708m4t1uRvFzK
bW2hwlvZCA8AW9QlEKz09Sggz7b6NIYFDSvtZFoGXL9glA0cfjPoNaWTbbHzFye08th8Ip0SRmMh
rqdW39E9B2vtbyOdhY0w8nOBIvq/vKHjaXy5Vkssiuk9FcaT++jYWSUhAAG+208Fy72zMZdLkohg
iJ8paIAww7DHTGuP6yjRMu61ay/DCxAOHVfZuwx3iM7QGS/hGDIBHgy7VpnsdrqQC1YFo4nQo9Ra
ugtGhkyr16UQtFicG9tNUP9ZgeP6ayt3f2UJp8nfBGd7GMcXMwj34WoUh98RGIgdRm1rGyZUn6cQ
Sa+eqm/V0xIEn2tRkz2c78T0B85HVD2Ejf2pyI9U15Q14xnpcGXkIxWDktwNFwgy/lgbHPagmgnc
rUUF8em0YAMjbrhG/99aNAnSMDSpGVga8S7WoZ7zNf99c9LCJMSG0otp0UXXCgbMVbxRmad96F7y
yZdSoyKQ9QLMVODGl+BJzlLfT7O2gd71UdzsIBll39KG0gIOaaN1xNdzT3542ulFY1YgFSBDKi4M
3R9+CiAjZ+rl8rCgisH/55SNKOAAKEDENoUfDIVNXP9pjTLev9wmZ0Njv9SLVH8bEmQ6890gFAfA
zV1ugigDRkVV+DQQNj5LbQnox+GbrOq3y+uMsSFn4pXXKs+AIHy6NR8ObvdfwheKdGNNiTC5oJ0k
w+tSqD5ij98jGAcw1BJfwtq1RRgI9PVffu7M4Jl0WGtR1Zr4CpFUjeZfUXhaoQVuP5tRiB0DZClb
XTAqwaM/0K3ChkXu0RXm5TfuuSVsC7oLYebY1XpNe9apAtTSf/Dxb7Lsa2Li01o/LAr4MmfbZIZr
ETu9NJIb+LGrR/YDOP59LPiYQf4zvlq7BMiW6T2p5pk1EqC8rWguAUEsBOsqbQzk9AucaKJvEk98
OgPVRAmKQP8/rH0/qKqpIfoCiAizRLgefGf3a0MorHzzNDlB9WHRWgQSSkdQh41Sywf+iBaR+VxA
n9/Zlc2tJDTuNfTJi6Dbt/wjlpY0ZQfyq9XPGzmjh+Re/ZtbAUvbmyqw4qzNZbwXnOSFgkMnwIMY
vrZlep67W/jf7NHoqCPv3I3HXaqePBjZEQMd6uIuj1LXQxkHJrH432TCF7g5q2ppllQB1aFSJpOQ
mudVJxbDdWMGCYYiZxhG8M+uLDkWJM7yvaybDNKIYnDu+VZgYEZT+Dse9/P0lG+NIHF65gD6skby
HI/NBtT+lyoHjyrd/C01aH8E2/Yr3Yi3N/4pF4Ey0KZAicSnxJr5HSAHXbiGHwAcAe7KISJLRBEl
l0MLnRU1DGHkUZIPfT/pjBzZLpbRD4386GKrNemZwsEZv7WWkDA2MkUF5r2zZd12D8YvJCsFe9sh
AVo6b4RDvEoX1GJYPJ77F0lCG4Ellqc9U4jZ4ex2WZIC3HFPR8TmXgD3wvLezv1vN3b4VgZ6v209
8iWIrX5ErcS+AiCQu29gi2j4A4moPE7xXWKdmVMxSh3mOUVRn1cjGR/gYaE3Of5sikxk+OxZOlOC
3vJ+p417XP/8YKpGa7Ds0ZYrsxF3TZ/gHnRCa/CS+1Rkwn0xzJ7EybriaV6QpCvoLgzWc0xpnL5K
YzI/GeRLN/Tizfiw2ZDSF5g6JbqkceeXuXg3DsZxWiUQBlAx3aA5fJTAbCwsLDtXu/kdqxsLg5Ab
evHOU21t0BO3GLNu7RD+dHl3k8fq27iY76JDZMRkFerh2gl5KNTydXDScRbNYYQ52GnxKttrE6WR
lf4MmNhCIV9ssdkfRJRMPTv5WphH1FdXBvnINt+zQDd9W2DeqfgdGmFg+8ipWPV+/cjRL7x4/30v
6b19zLSpsYjTjky6cfdWJtBupJqI03DuH6r9IBSZnui6YDy2wQ0L0T5ZWNqYGAleuLgdzequ7KSr
DzYyWHmcyXH9EyhnNMpl7LwGsedalfHzqlf6O6TZh96mSetBTsEzhGF0O0y2Cc06Q4l4oVM4KkMn
kWOFJ5w6W2/qhADsLH229N9095b+DxhdZ+u2+CVUKQy+F2QlUBwZEMvAvWcdhw47A2n2I0yMWavR
cV6aYePezeLlktvpXFzFLcKFMWLPAubsmiWI2YF/tCYNyOSqq5702LXldFulM7iglk5K1miMsFcI
JaVZIK2JFMpJk2NIKQQq32hJxwGvFam5C818L8NTRx5Ad2M/zg86ZAqnCzkmeLn2c0/zADhfEbij
B3v7RR6d0jSVNpV5djtmOEiftQE7sNAvKSkzUF3U8C3y+FMfGPLpZ8Fd0o+nZ3eV7QQXE2u9Muyh
5t92sA2LvDHxEkytWSMBNgPDcdLQojYiBzERywY9nSBfIqr6McThB79mecixtVDwGKSxPAwW4zJe
40ozrnmF2DccEYqWwm8A4vmOBrLBL+v6oZANiyRiKrjd2o5AwZehKKsFfhHgaKLjwoyYn0DFPoGc
lHmAajEdWqHZ/bKonqiB3L23w75C+MUn00uoDK2NKrGCPK8Sds3opYuM5NIfZ67ZpZjbAzJqLZBw
mFZwkZzpkq40We1omaOt1acQG5Cr2pV0bayismldMR6Q085yd0lF3f5Wkiq9Y0ZtEjAkIwh8nmXX
zkj/2exiXPEWAvLp/oec7XDMc/63fFmpGknyG1mzONj0YaDIz2hrMyvu0cTNhvQ7xiqxTgeEV4uI
CfPR6VXc+FNGzcOxavv+RN5WZ1SxJPU=
`pragma protect end_protected
